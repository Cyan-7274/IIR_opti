
module opti_top ( clk, rst_n, data_in, valid_in, data_out, valid_out );
  input [15:0] data_in;
  output [15:0] data_out;
  input clk, rst_n, valid_in;
  output valid_out;
  wire   \sos_data[1][15] , \sos_data[1][14] , \sos_data[1][13] ,
         \sos_data[1][12] , \sos_data[1][11] , \sos_data[1][10] ,
         \sos_data[1][9] , \sos_data[1][8] , \sos_data[1][7] ,
         \sos_data[1][6] , \sos_data[1][5] , \sos_data[1][4] ,
         \sos_data[1][3] , \sos_data[1][2] , \sos_data[1][1] ,
         \sos_data[1][0] , \sos_data[2][15] , \sos_data[2][14] ,
         \sos_data[2][13] , \sos_data[2][12] , \sos_data[2][11] ,
         \sos_data[2][10] , \sos_data[2][9] , \sos_data[2][8] ,
         \sos_data[2][7] , \sos_data[2][6] , \sos_data[2][5] ,
         \sos_data[2][4] , \sos_data[2][3] , \sos_data[2][2] ,
         \sos_data[2][1] , \sos_data[2][0] , \sos_data[3][15] ,
         \sos_data[3][14] , \sos_data[3][13] , \sos_data[3][12] ,
         \sos_data[3][11] , \sos_data[3][10] , \sos_data[3][9] ,
         \sos_data[3][8] , \sos_data[3][7] , \sos_data[3][6] ,
         \sos_data[3][5] , \sos_data[3][4] , \sos_data[3][3] ,
         \sos_data[3][2] , \sos_data[3][1] , \sos_data[3][0] ,
         \sos_data[4][15] , \sos_data[4][14] , \sos_data[4][13] ,
         \sos_data[4][12] , \sos_data[4][11] , \sos_data[4][10] ,
         \sos_data[4][9] , \sos_data[4][8] , \sos_data[4][7] ,
         \sos_data[4][6] , \sos_data[4][5] , \sos_data[4][4] ,
         \sos_data[4][3] , \sos_data[4][2] , \sos_data[4][1] ,
         \sos_data[4][0] , net199029, net199030, net199031, net199032,
         net199033, net199034, net199035, net199036, net199037, net199038,
         net199039, net199040, net199041, net199042, net199043, net199044,
         net199045, net199046, net199047, net199048, net199049, net199050,
         net199051, net199052, net199053, net199054, net199055, net199056,
         net199057, net199058, net199059, net199060, net199061, net199062,
         net199063, net199064, net199065, net199066, net199067, net199068,
         net199069, net199070, net199071, net199072, net199073, net199074,
         net199075, net199076, net199077, net199078, net199079, net199080,
         net199081, net199082, net199083, net199084, net199085, net199086,
         net199087, net199088, net199089, net199090, net199091, net199092,
         net199093, net199094, net199095, net199096, net199097, net199098,
         net199099, net199100, net199101, net199102, net199103, net199104,
         net199105, net199106, net199107, net199108, net199109, net199110,
         net199111, net199112, net199113, net199114, net199115, net199116,
         net199117, net199118, net199119, net199120, net199121, net199122,
         net199123, net199124, net199125, net199126, net199127, net199128,
         net199129, net199130, net199131, net199132, net199133, net199134,
         net199135, net199136, net199137, net199138, net199139, net199140,
         net199141, net199142, net199143, net199144, net199145, net199146,
         net199147, net199148, net199149, net199150, net199151, net199152,
         net199153, net199154, net199155, net199156, net199157, net199158,
         net199159, net199160, net199161, net199162, net199163, net199164,
         net199165, net199166, net199167, net199168, net199169, net199170,
         net199171, net199172, net199173, net199174, net199175, net199176,
         net199177, net199178, net199179, net199180, net199181, net199182,
         net199183, net199184, net199185, net199186, net199187, net199188,
         net199189, net199190, net199191, net199192, net199193, net199194,
         net199195, net199196, net199197, net199198, net199199, net199200,
         net199201, net199202, net199203, net199204, net199205, net199206,
         net199207, net199208, net199209, net199210, net199211, net199212,
         net199213, net199214, net199215, net199216, net199217, net199218,
         net199219, net199220, net199221, net199222, net199223, net199224,
         net199225, net199226, net199227, net199228, net199229, net199230,
         net199231, net199232, net199233, net199234, net199235, net199236,
         net199237, net199238, net199239, net199240, net199241, net199242,
         net199243, net199244, net199245, net199246, net199247, net199248,
         net199249, net199250, net199251, net199252, net199253, net199254,
         net199255, net199256, net199257, net199258, net199259, net199260,
         net199261, net199262, net199263, net199264, net199265, net199266,
         net199267, net199268, net199269, net199270, net199271, net199272,
         net199273, net199274, net199275, net199276, net199277, net199278,
         net199279, net199280, net199281, net199282, net199283, net199284,
         net199285, net199286, net199287, net199288, net199289, net199290,
         net199291, net199292, net199293, net199294, net199295, net199296,
         net199297, net199298, net199299, net199300, net199301, net199302,
         net199303, net199304, net199305, net199306, net199307, net199308,
         net199309, net199310, net199311, net199312, net199313, net199314,
         net199315, net199316, net199317, net199318, net199319, net199320,
         net199321, net199322, net199323, net199324, net199325, net199326,
         net199327, net199328, net199329, net199330, net199331, net199332,
         net199333, net199334, net199335, net199336, net199337, net199338,
         net199339, net199340, net199341, net199342, net199343, net199344,
         net199345, net199346, net199347, net199348, net199349, net199350,
         net199351, net199352, net199353, net199354, net199355, net199356,
         net199357, net199358, net199359, net199360, net199361, net199362,
         net199363, net199364, net199365, net199366, net199367, net199368,
         net199369, net199370, net199371, net199372, net199373, net199374,
         net199375, net199376, net199377, net199378, net199379, net199380,
         net199381, net199382, net199383, net199384, net199385, net199386,
         net199387, net199388, net199389, net199390, net199391, net199392,
         net199393, net199394, net199395, net199396, net199397, net199398,
         net199399, net199400, net199401, net199402, net199403, net199404,
         net199405, net199406, net199407, net199408, net199409, net199410,
         net199411, net199412, net199413, net199414, net199415, net199416,
         net199417, net199418, net199419, net199420, net199421, net199422,
         net199423, net199424, net199425, net199426, net199427, net199428;
  wire   [1:4] sos_valid;

  opti_sos_0 \SOS_CHAIN[0].u_sos  ( .clk(clk), .rst_n(rst_n), .data_in(data_in), .valid_in(valid_in), .b0({net199349, net199350, net199351, net199352, 
        net199353, net199354, net199355, net199356, net199357, net199358, 
        net199359, net199360, net199361, net199362, net199363, net199364}), 
        .b1({net199365, net199366, net199367, net199368, net199369, net199370, 
        net199371, net199372, net199373, net199374, net199375, net199376, 
        net199377, net199378, net199379, net199380}), .b2({net199381, 
        net199382, net199383, net199384, net199385, net199386, net199387, 
        net199388, net199389, net199390, net199391, net199392, net199393, 
        net199394, net199395, net199396}), .a1({net199397, net199398, 
        net199399, net199400, net199401, net199402, net199403, net199404, 
        net199405, net199406, net199407, net199408, net199409, net199410, 
        net199411, net199412}), .a2({net199413, net199414, net199415, 
        net199416, net199417, net199418, net199419, net199420, net199421, 
        net199422, net199423, net199424, net199425, net199426, net199427, 
        net199428}), .data_out({\sos_data[1][15] , \sos_data[1][14] , 
        \sos_data[1][13] , \sos_data[1][12] , \sos_data[1][11] , 
        \sos_data[1][10] , \sos_data[1][9] , \sos_data[1][8] , 
        \sos_data[1][7] , \sos_data[1][6] , \sos_data[1][5] , \sos_data[1][4] , 
        \sos_data[1][3] , \sos_data[1][2] , \sos_data[1][1] , \sos_data[1][0] }), .valid_out(sos_valid[1]) );
  opti_sos_4 \SOS_CHAIN[1].u_sos  ( .clk(clk), .rst_n(rst_n), .data_in({
        \sos_data[1][15] , \sos_data[1][14] , \sos_data[1][13] , 
        \sos_data[1][12] , \sos_data[1][11] , \sos_data[1][10] , 
        \sos_data[1][9] , \sos_data[1][8] , \sos_data[1][7] , \sos_data[1][6] , 
        \sos_data[1][5] , \sos_data[1][4] , \sos_data[1][3] , \sos_data[1][2] , 
        \sos_data[1][1] , \sos_data[1][0] }), .valid_in(sos_valid[1]), .b0({
        net199269, net199270, net199271, net199272, net199273, net199274, 
        net199275, net199276, net199277, net199278, net199279, net199280, 
        net199281, net199282, net199283, net199284}), .b1({net199285, 
        net199286, net199287, net199288, net199289, net199290, net199291, 
        net199292, net199293, net199294, net199295, net199296, net199297, 
        net199298, net199299, net199300}), .b2({net199301, net199302, 
        net199303, net199304, net199305, net199306, net199307, net199308, 
        net199309, net199310, net199311, net199312, net199313, net199314, 
        net199315, net199316}), .a1({net199317, net199318, net199319, 
        net199320, net199321, net199322, net199323, net199324, net199325, 
        net199326, net199327, net199328, net199329, net199330, net199331, 
        net199332}), .a2({net199333, net199334, net199335, net199336, 
        net199337, net199338, net199339, net199340, net199341, net199342, 
        net199343, net199344, net199345, net199346, net199347, net199348}), 
        .data_out({\sos_data[2][15] , \sos_data[2][14] , \sos_data[2][13] , 
        \sos_data[2][12] , \sos_data[2][11] , \sos_data[2][10] , 
        \sos_data[2][9] , \sos_data[2][8] , \sos_data[2][7] , \sos_data[2][6] , 
        \sos_data[2][5] , \sos_data[2][4] , \sos_data[2][3] , \sos_data[2][2] , 
        \sos_data[2][1] , \sos_data[2][0] }), .valid_out(sos_valid[2]) );
  opti_sos_3 \SOS_CHAIN[2].u_sos  ( .clk(clk), .rst_n(rst_n), .data_in({
        \sos_data[2][15] , \sos_data[2][14] , \sos_data[2][13] , 
        \sos_data[2][12] , \sos_data[2][11] , \sos_data[2][10] , 
        \sos_data[2][9] , \sos_data[2][8] , \sos_data[2][7] , \sos_data[2][6] , 
        \sos_data[2][5] , \sos_data[2][4] , \sos_data[2][3] , \sos_data[2][2] , 
        \sos_data[2][1] , \sos_data[2][0] }), .valid_in(sos_valid[2]), .b0({
        net199189, net199190, net199191, net199192, net199193, net199194, 
        net199195, net199196, net199197, net199198, net199199, net199200, 
        net199201, net199202, net199203, net199204}), .b1({net199205, 
        net199206, net199207, net199208, net199209, net199210, net199211, 
        net199212, net199213, net199214, net199215, net199216, net199217, 
        net199218, net199219, net199220}), .b2({net199221, net199222, 
        net199223, net199224, net199225, net199226, net199227, net199228, 
        net199229, net199230, net199231, net199232, net199233, net199234, 
        net199235, net199236}), .a1({net199237, net199238, net199239, 
        net199240, net199241, net199242, net199243, net199244, net199245, 
        net199246, net199247, net199248, net199249, net199250, net199251, 
        net199252}), .a2({net199253, net199254, net199255, net199256, 
        net199257, net199258, net199259, net199260, net199261, net199262, 
        net199263, net199264, net199265, net199266, net199267, net199268}), 
        .data_out({\sos_data[3][15] , \sos_data[3][14] , \sos_data[3][13] , 
        \sos_data[3][12] , \sos_data[3][11] , \sos_data[3][10] , 
        \sos_data[3][9] , \sos_data[3][8] , \sos_data[3][7] , \sos_data[3][6] , 
        \sos_data[3][5] , \sos_data[3][4] , \sos_data[3][3] , \sos_data[3][2] , 
        \sos_data[3][1] , \sos_data[3][0] }), .valid_out(sos_valid[3]) );
  opti_sos_2 \SOS_CHAIN[3].u_sos  ( .clk(clk), .rst_n(rst_n), .data_in({
        \sos_data[3][15] , \sos_data[3][14] , \sos_data[3][13] , 
        \sos_data[3][12] , \sos_data[3][11] , \sos_data[3][10] , 
        \sos_data[3][9] , \sos_data[3][8] , \sos_data[3][7] , \sos_data[3][6] , 
        \sos_data[3][5] , \sos_data[3][4] , \sos_data[3][3] , \sos_data[3][2] , 
        \sos_data[3][1] , \sos_data[3][0] }), .valid_in(sos_valid[3]), .b0({
        net199109, net199110, net199111, net199112, net199113, net199114, 
        net199115, net199116, net199117, net199118, net199119, net199120, 
        net199121, net199122, net199123, net199124}), .b1({net199125, 
        net199126, net199127, net199128, net199129, net199130, net199131, 
        net199132, net199133, net199134, net199135, net199136, net199137, 
        net199138, net199139, net199140}), .b2({net199141, net199142, 
        net199143, net199144, net199145, net199146, net199147, net199148, 
        net199149, net199150, net199151, net199152, net199153, net199154, 
        net199155, net199156}), .a1({net199157, net199158, net199159, 
        net199160, net199161, net199162, net199163, net199164, net199165, 
        net199166, net199167, net199168, net199169, net199170, net199171, 
        net199172}), .a2({net199173, net199174, net199175, net199176, 
        net199177, net199178, net199179, net199180, net199181, net199182, 
        net199183, net199184, net199185, net199186, net199187, net199188}), 
        .data_out({\sos_data[4][15] , \sos_data[4][14] , \sos_data[4][13] , 
        \sos_data[4][12] , \sos_data[4][11] , \sos_data[4][10] , 
        \sos_data[4][9] , \sos_data[4][8] , \sos_data[4][7] , \sos_data[4][6] , 
        \sos_data[4][5] , \sos_data[4][4] , \sos_data[4][3] , \sos_data[4][2] , 
        \sos_data[4][1] , \sos_data[4][0] }), .valid_out(sos_valid[4]) );
  opti_sos_1 \SOS_CHAIN[4].u_sos  ( .clk(clk), .rst_n(rst_n), .data_in({
        \sos_data[4][15] , \sos_data[4][14] , \sos_data[4][13] , 
        \sos_data[4][12] , \sos_data[4][11] , \sos_data[4][10] , 
        \sos_data[4][9] , \sos_data[4][8] , \sos_data[4][7] , \sos_data[4][6] , 
        \sos_data[4][5] , \sos_data[4][4] , \sos_data[4][3] , \sos_data[4][2] , 
        \sos_data[4][1] , \sos_data[4][0] }), .valid_in(sos_valid[4]), .b0({
        net199029, net199030, net199031, net199032, net199033, net199034, 
        net199035, net199036, net199037, net199038, net199039, net199040, 
        net199041, net199042, net199043, net199044}), .b1({net199045, 
        net199046, net199047, net199048, net199049, net199050, net199051, 
        net199052, net199053, net199054, net199055, net199056, net199057, 
        net199058, net199059, net199060}), .b2({net199061, net199062, 
        net199063, net199064, net199065, net199066, net199067, net199068, 
        net199069, net199070, net199071, net199072, net199073, net199074, 
        net199075, net199076}), .a1({net199077, net199078, net199079, 
        net199080, net199081, net199082, net199083, net199084, net199085, 
        net199086, net199087, net199088, net199089, net199090, net199091, 
        net199092}), .a2({net199093, net199094, net199095, net199096, 
        net199097, net199098, net199099, net199100, net199101, net199102, 
        net199103, net199104, net199105, net199106, net199107, net199108}), 
        .data_out(data_out), .valid_out(valid_out) );
endmodule


module opti_sos_4 ( clk, rst_n, data_in, valid_in, b0, b1, b2, a1, a2, 
        data_out, valid_out );
  input [15:0] data_in;
  input [15:0] b0;
  input [15:0] b1;
  input [15:0] b2;
  input [15:0] a1;
  input [15:0] a2;
  output [15:0] data_out;
  input clk, rst_n, valid_in;
  output valid_out;
  wire   valid_T1, valid_T3, valid_T2, \mul_b0/result_sat[15] ,
         \mul_b0/result_sat[14] , \mul_b0/result_sat[13] ,
         \mul_b0/result_sat[12] , \mul_b0/result_sat[11] ,
         \mul_b0/result_sat[10] , \mul_b0/result_sat[9] ,
         \mul_b0/result_sat[8] , \mul_b0/result_sat[7] ,
         \mul_b0/result_sat[6] , \mul_b0/result_sat[5] ,
         \mul_b0/result_sat[4] , \mul_b0/result_sat[3] ,
         \mul_b0/result_sat[2] , \mul_b0/result_sat[1] ,
         \mul_b0/result_sat[0] , \mul_b0/fa1_s2_r[33] , \mul_b0/fa1_s2_r[32] ,
         \mul_b0/fa1_s2_r[31] , \mul_b0/fa1_s2_r[30] , \mul_b0/fa1_s2_r[29] ,
         \mul_b0/fa1_s2_r[28] , \mul_b0/fa1_s2_r[27] , \mul_b0/fa1_s2_r[26] ,
         \mul_b0/fa1_s2_r[25] , \mul_b0/fa1_s2_r[24] , \mul_b0/fa1_s2_r[23] ,
         \mul_b0/fa1_s2_r[22] , \mul_b0/fa1_s2_r[21] , \mul_b0/fa1_s2_r[20] ,
         \mul_b0/fa1_s2_r[19] , \mul_b0/fa1_s2_r[18] , \mul_b0/fa1_s2_r[17] ,
         \mul_b0/fa1_s2_r[16] , \mul_b0/fa1_s2_r[15] , \mul_b0/fa1_s2_r[14] ,
         \mul_b0/fa1_s2_r[13] , \mul_b0/fa1_s2_r[12] , \mul_b0/fa1_s1_r[33] ,
         \mul_b0/fa1_s1_r[32] , \mul_b0/fa1_s1_r[31] , \mul_b0/fa1_s1_r[30] ,
         \mul_b0/fa1_s1_r[29] , \mul_b0/fa1_s1_r[28] , \mul_b0/fa1_s1_r[27] ,
         \mul_b0/fa1_s1_r[26] , \mul_b0/fa1_s1_r[25] , \mul_b0/fa1_s1_r[24] ,
         \mul_b0/fa1_s1_r[23] , \mul_b0/fa1_s1_r[22] , \mul_b0/fa1_s1_r[21] ,
         \mul_b0/fa1_s1_r[20] , \mul_b0/fa1_s1_r[19] , \mul_b0/fa1_s1_r[18] ,
         \mul_b0/fa1_s1_r[17] , \mul_b0/fa1_s1_r[16] , \mul_b0/fa1_s1_r[15] ,
         \mul_b0/fa1_s1_r[14] , \mul_b0/fa1_s1_r[13] , \mul_b0/fa1_s1_r[12] ,
         \mul_b0/fa1_s1_r[11] , \mul_b0/fa1_s1_r[10] , \mul_b0/fa1_s1_r[9] ,
         \mul_b0/fa1_s1_r[8] , \mul_b0/fa1_c0_r[20] , \mul_b0/fa1_c0_r[19] ,
         \mul_b0/fa1_c0_r[18] , \mul_b0/fa1_c0_r[17] , \mul_b0/fa1_c0_r[16] ,
         \mul_b0/fa1_c0_r[15] , \mul_b0/fa1_c0_r[14] , \mul_b0/fa1_c0_r[13] ,
         \mul_b0/fa1_c0_r[12] , \mul_b0/fa1_c0_r[11] , \mul_b0/fa1_c0_r[10] ,
         \mul_b0/fa1_c0_r[9] , \mul_b0/fa1_c0_r[8] , \mul_b0/fa1_c0_r[7] ,
         \mul_b0/fa1_c0_r[6] , \mul_b0/fa1_c0_r[5] , \mul_b0/fa1_s0_r[33] ,
         \mul_b0/fa1_s0_r[32] , \mul_b0/fa1_s0_r[31] , \mul_b0/fa1_s0_r[30] ,
         \mul_b0/fa1_s0_r[29] , \mul_b0/fa1_s0_r[28] , \mul_b0/fa1_s0_r[27] ,
         \mul_b0/fa1_s0_r[26] , \mul_b0/fa1_s0_r[25] , \mul_b0/fa1_s0_r[24] ,
         \mul_b0/fa1_s0_r[23] , \mul_b0/fa1_s0_r[22] , \mul_b0/fa1_s0_r[21] ,
         \mul_b0/fa1_s0_r[20] , \mul_b0/fa1_s0_r[19] , \mul_b0/fa1_s0_r[18] ,
         \mul_b0/fa1_s0_r[17] , \mul_b0/fa1_s0_r[16] , \mul_b0/fa1_s0_r[15] ,
         \mul_b0/fa1_s0_r[14] , \mul_b0/fa1_s0_r[13] , \mul_b0/fa1_s0_r[12] ,
         \mul_b0/fa1_s0_r[11] , \mul_b0/fa1_s0_r[10] , \mul_b0/fa1_s0_r[9] ,
         \mul_b0/fa1_s0_r[8] , \mul_b0/fa1_s0_r[7] , \mul_b0/fa1_s0_r[6] ,
         \mul_b0/fa1_c0[20] , \mul_b0/fa1_c0[19] , \mul_b0/fa1_c0[18] ,
         \mul_b0/fa1_c0[17] , \mul_b0/fa1_c0[16] , \mul_b0/fa1_c0[15] ,
         \mul_b0/fa1_c0[14] , \mul_b0/fa1_c0[13] , \mul_b0/fa1_c0[12] ,
         \mul_b0/fa1_c0[11] , \mul_b0/fa1_c0[10] , \mul_b0/fa1_c0[9] ,
         \mul_b0/fa1_c0[8] , \mul_b0/fa1_c0[7] , \mul_b0/fa1_c0[6] ,
         \mul_b0/fa1_c0[5] , \mul_b0/fa1_s0[30] , \mul_b0/fa1_s0[20] ,
         \mul_b0/fa1_s0[19] , \mul_b0/fa1_s0[18] , \mul_b0/fa1_s0[17] ,
         \mul_b0/fa1_s0[16] , \mul_b0/fa1_s0[15] , \mul_b0/fa1_s0[14] ,
         \mul_b0/fa1_s0[13] , \mul_b0/fa1_s0[12] , \mul_b0/fa1_s0[11] ,
         \mul_b0/fa1_s0[10] , \mul_b0/fa1_s0[9] , \mul_b0/fa1_s0[8] ,
         \mul_b0/fa1_s0[7] , \mul_b0/fa1_s0[6] , \mul_b1/result_sat[15] ,
         \mul_b1/result_sat[14] , \mul_b1/result_sat[13] ,
         \mul_b1/result_sat[12] , \mul_b1/result_sat[11] ,
         \mul_b1/result_sat[10] , \mul_b1/result_sat[9] ,
         \mul_b1/result_sat[8] , \mul_b1/result_sat[7] ,
         \mul_b1/result_sat[6] , \mul_b1/result_sat[5] ,
         \mul_b1/result_sat[4] , \mul_b1/result_sat[3] ,
         \mul_b1/result_sat[2] , \mul_b1/result_sat[1] ,
         \mul_b1/result_sat[0] , \mul_b1/fa1_c2_r[28] , \mul_b1/fa1_c2_r[27] ,
         \mul_b1/fa1_c2_r[26] , \mul_b1/fa1_c2_r[25] , \mul_b1/fa1_c2_r[24] ,
         \mul_b1/fa1_c2_r[23] , \mul_b1/fa1_c2_r[22] , \mul_b1/fa1_c2_r[21] ,
         \mul_b1/fa1_c2_r[20] , \mul_b1/fa1_c2_r[19] , \mul_b1/fa1_c2_r[18] ,
         \mul_b1/fa1_c2_r[17] , \mul_b1/fa1_c2_r[16] , \mul_b1/fa1_c2_r[15] ,
         \mul_b1/fa1_c2_r[14] , \mul_b1/fa1_s2_r[33] , \mul_b1/fa1_s2_r[32] ,
         \mul_b1/fa1_s2_r[31] , \mul_b1/fa1_s2_r[30] , \mul_b1/fa1_s2_r[29] ,
         \mul_b1/fa1_s2_r[28] , \mul_b1/fa1_s2_r[27] , \mul_b1/fa1_s2_r[26] ,
         \mul_b1/fa1_s2_r[25] , \mul_b1/fa1_s2_r[24] , \mul_b1/fa1_s2_r[23] ,
         \mul_b1/fa1_s2_r[22] , \mul_b1/fa1_s2_r[21] , \mul_b1/fa1_s2_r[20] ,
         \mul_b1/fa1_s2_r[19] , \mul_b1/fa1_s2_r[18] , \mul_b1/fa1_s2_r[17] ,
         \mul_b1/fa1_s2_r[16] , \mul_b1/fa1_s2_r[15] , \mul_b1/fa1_s2_r[14] ,
         \mul_b1/fa1_s2_r[13] , \mul_b1/fa1_c1_r[32] , \mul_b1/fa1_c1_r[31] ,
         \mul_b1/fa1_c1_r[30] , \mul_b1/fa1_c1_r[29] , \mul_b1/fa1_c1_r[28] ,
         \mul_b1/fa1_c1_r[27] , \mul_b1/fa1_c1_r[26] , \mul_b1/fa1_c1_r[25] ,
         \mul_b1/fa1_c1_r[24] , \mul_b1/fa1_c1_r[23] , \mul_b1/fa1_c1_r[22] ,
         \mul_b1/fa1_c1_r[21] , \mul_b1/fa1_c1_r[20] , \mul_b1/fa1_c1_r[19] ,
         \mul_b1/fa1_c1_r[18] , \mul_b1/fa1_c1_r[17] , \mul_b1/fa1_c1_r[16] ,
         \mul_b1/fa1_c1_r[15] , \mul_b1/fa1_c1_r[14] , \mul_b1/fa1_c1_r[13] ,
         \mul_b1/fa1_c1_r[12] , \mul_b1/fa1_c1_r[11] , \mul_b1/fa1_c1_r[10] ,
         \mul_b1/fa1_c1_r[9] , \mul_b1/fa1_c1_r[8] , \mul_b1/fa1_s1_r[33] ,
         \mul_b1/fa1_s1_r[32] , \mul_b1/fa1_s1_r[31] , \mul_b1/fa1_s1_r[30] ,
         \mul_b1/fa1_s1_r[29] , \mul_b1/fa1_s1_r[28] , \mul_b1/fa1_s1_r[27] ,
         \mul_b1/fa1_s1_r[26] , \mul_b1/fa1_s1_r[25] , \mul_b1/fa1_s1_r[24] ,
         \mul_b1/fa1_s1_r[23] , \mul_b1/fa1_s1_r[22] , \mul_b1/fa1_s1_r[21] ,
         \mul_b1/fa1_s1_r[20] , \mul_b1/fa1_s1_r[19] , \mul_b1/fa1_s1_r[18] ,
         \mul_b1/fa1_s1_r[17] , \mul_b1/fa1_s1_r[16] , \mul_b1/fa1_s1_r[15] ,
         \mul_b1/fa1_s1_r[14] , \mul_b1/fa1_s1_r[13] , \mul_b1/fa1_s1_r[12] ,
         \mul_b1/fa1_s1_r[11] , \mul_b1/fa1_s1_r[10] , \mul_b1/fa1_s1_r[9] ,
         \mul_b1/fa1_s1_r[8] , \mul_b1/fa1_s1_r[7] , \mul_b1/fa1_s1_r[6] ,
         \mul_b1/fa1_c0_r[32] , \mul_b1/fa1_c0_r[31] , \mul_b1/fa1_c0_r[30] ,
         \mul_b1/fa1_c0_r[29] , \mul_b1/fa1_c0_r[28] , \mul_b1/fa1_c0_r[27] ,
         \mul_b1/fa1_c0_r[26] , \mul_b1/fa1_c0_r[25] , \mul_b1/fa1_c0_r[24] ,
         \mul_b1/fa1_c0_r[23] , \mul_b1/fa1_c0_r[22] , \mul_b1/fa1_c0_r[21] ,
         \mul_b1/fa1_c0_r[20] , \mul_b1/fa1_c0_r[19] , \mul_b1/fa1_c0_r[18] ,
         \mul_b1/fa1_c0_r[17] , \mul_b1/fa1_c0_r[16] , \mul_b1/fa1_c0_r[15] ,
         \mul_b1/fa1_c0_r[14] , \mul_b1/fa1_c0_r[13] , \mul_b1/fa1_c0_r[12] ,
         \mul_b1/fa1_c0_r[11] , \mul_b1/fa1_c0_r[10] , \mul_b1/fa1_c0_r[9] ,
         \mul_b1/fa1_c0_r[8] , \mul_b1/fa1_c0_r[7] , \mul_b1/fa1_c0_r[6] ,
         \mul_b1/fa1_c0_r[5] , \mul_b1/fa1_c0_r[4] , \mul_b1/fa1_c0_r[3] ,
         \mul_b1/fa1_c0_r[2] , \mul_b1/fa1_s0_r[33] , \mul_b1/fa1_s0_r[32] ,
         \mul_b1/fa1_s0_r[31] , \mul_b1/fa1_s0_r[30] , \mul_b1/fa1_s0_r[29] ,
         \mul_b1/fa1_s0_r[28] , \mul_b1/fa1_s0_r[27] , \mul_b1/fa1_s0_r[26] ,
         \mul_b1/fa1_s0_r[25] , \mul_b1/fa1_s0_r[24] , \mul_b1/fa1_s0_r[23] ,
         \mul_b1/fa1_s0_r[22] , \mul_b1/fa1_s0_r[21] , \mul_b1/fa1_s0_r[20] ,
         \mul_b1/fa1_s0_r[19] , \mul_b1/fa1_s0_r[18] , \mul_b1/fa1_s0_r[17] ,
         \mul_b1/fa1_s0_r[16] , \mul_b1/fa1_s0_r[15] , \mul_b1/fa1_s0_r[14] ,
         \mul_b1/fa1_s0_r[13] , \mul_b1/fa1_s0_r[12] , \mul_b1/fa1_s0_r[11] ,
         \mul_b1/fa1_s0_r[10] , \mul_b1/fa1_s0_r[9] , \mul_b1/fa1_s0_r[8] ,
         \mul_b1/fa1_s0_r[7] , \mul_b1/fa1_s0_r[6] , \mul_b1/fa1_s0_r[5] ,
         \mul_b1/fa1_s0_r[4] , \mul_b1/fa1_s0_r[3] , \mul_b1/fa1_c2[28] ,
         \mul_b1/fa1_c2[27] , \mul_b1/fa1_c2[26] , \mul_b1/fa1_c2[25] ,
         \mul_b1/fa1_c2[24] , \mul_b1/fa1_c2[23] , \mul_b1/fa1_c2[22] ,
         \mul_b1/fa1_c2[21] , \mul_b1/fa1_c2[20] , \mul_b1/fa1_c2[19] ,
         \mul_b1/fa1_c2[18] , \mul_b1/fa1_c2[17] , \mul_b1/fa1_c2[16] ,
         \mul_b1/fa1_c2[15] , \mul_b1/fa1_c2[14] , \mul_b1/fa1_s2[29] ,
         \mul_b1/fa1_s2[28] , \mul_b1/fa1_s2[27] , \mul_b1/fa1_s2[26] ,
         \mul_b1/fa1_s2[25] , \mul_b1/fa1_s2[24] , \mul_b1/fa1_s2[23] ,
         \mul_b1/fa1_s2[22] , \mul_b1/fa1_s2[21] , \mul_b1/fa1_s2[20] ,
         \mul_b1/fa1_s2[19] , \mul_b1/fa1_s2[18] , \mul_b1/fa1_s2[17] ,
         \mul_b1/fa1_s2[16] , \mul_b1/fa1_s2[15] , \mul_b1/fa1_s2[14] ,
         \mul_b1/fa1_c1[22] , \mul_b1/fa1_c1[21] , \mul_b1/fa1_c1[20] ,
         \mul_b1/fa1_c1[19] , \mul_b1/fa1_c1[18] , \mul_b1/fa1_c1[17] ,
         \mul_b1/fa1_c1[16] , \mul_b1/fa1_c1[15] , \mul_b1/fa1_c1[14] ,
         \mul_b1/fa1_c1[13] , \mul_b1/fa1_c1[12] , \mul_b1/fa1_c1[11] ,
         \mul_b1/fa1_c1[10] , \mul_b1/fa1_c1[9] , \mul_b1/fa1_c1[8] ,
         \mul_b1/fa1_s1[25] , \mul_b1/fa1_s1[24] , \mul_b1/fa1_s1[23] ,
         \mul_b1/fa1_s1[22] , \mul_b1/fa1_s1[21] , \mul_b1/fa1_s1[20] ,
         \mul_b1/fa1_s1[19] , \mul_b1/fa1_s1[18] , \mul_b1/fa1_s1[17] ,
         \mul_b1/fa1_s1[16] , \mul_b1/fa1_s1[15] , \mul_b1/fa1_s1[14] ,
         \mul_b1/fa1_s1[13] , \mul_b1/fa1_s1[12] , \mul_b1/fa1_s1[11] ,
         \mul_b1/fa1_s1[10] , \mul_b1/fa1_s1[9] , \mul_b1/fa1_s1[8] ,
         \mul_b1/fa1_s1[7] , \mul_b1/fa1_c0[16] , \mul_b1/fa1_c0[15] ,
         \mul_b1/fa1_c0[14] , \mul_b1/fa1_c0[13] , \mul_b1/fa1_c0[12] ,
         \mul_b1/fa1_c0[11] , \mul_b1/fa1_c0[10] , \mul_b1/fa1_c0[9] ,
         \mul_b1/fa1_c0[8] , \mul_b1/fa1_c0[7] , \mul_b1/fa1_c0[6] ,
         \mul_b1/fa1_c0[5] , \mul_b1/fa1_s0[16] , \mul_b1/fa1_s0[15] ,
         \mul_b1/fa1_s0[14] , \mul_b1/fa1_s0[13] , \mul_b1/fa1_s0[12] ,
         \mul_b1/fa1_s0[11] , \mul_b1/fa1_s0[10] , \mul_b1/fa1_s0[9] ,
         \mul_b1/fa1_s0[8] , \mul_b1/fa1_s0[7] , \mul_b1/fa1_s0[6] ,
         \mul_b1/fa1_s0[5] , \mul_b1/fa1_s0[4] , \mul_b1/fa1_s0[3] ,
         \mul_b2/result_sat[15] , \mul_b2/result_sat[14] ,
         \mul_b2/result_sat[13] , \mul_b2/result_sat[12] ,
         \mul_b2/result_sat[11] , \mul_b2/result_sat[10] ,
         \mul_b2/result_sat[9] , \mul_b2/result_sat[8] ,
         \mul_b2/result_sat[7] , \mul_b2/result_sat[6] ,
         \mul_b2/result_sat[5] , \mul_b2/result_sat[4] ,
         \mul_b2/result_sat[3] , \mul_b2/result_sat[2] ,
         \mul_b2/result_sat[1] , \mul_b2/result_sat[0] , \mul_b2/fa1_s2_r[33] ,
         \mul_b2/fa1_s2_r[32] , \mul_b2/fa1_s2_r[31] , \mul_b2/fa1_s2_r[30] ,
         \mul_b2/fa1_s2_r[29] , \mul_b2/fa1_s2_r[28] , \mul_b2/fa1_s2_r[27] ,
         \mul_b2/fa1_s2_r[26] , \mul_b2/fa1_s2_r[25] , \mul_b2/fa1_s2_r[24] ,
         \mul_b2/fa1_s2_r[23] , \mul_b2/fa1_s2_r[22] , \mul_b2/fa1_s2_r[21] ,
         \mul_b2/fa1_s2_r[20] , \mul_b2/fa1_s2_r[19] , \mul_b2/fa1_s2_r[18] ,
         \mul_b2/fa1_s2_r[17] , \mul_b2/fa1_s2_r[16] , \mul_b2/fa1_s2_r[15] ,
         \mul_b2/fa1_s2_r[14] , \mul_b2/fa1_s2_r[13] , \mul_b2/fa1_s2_r[12] ,
         \mul_b2/fa1_c1_r[23] , \mul_b2/fa1_c1_r[22] , \mul_b2/fa1_c1_r[21] ,
         \mul_b2/fa1_c1_r[20] , \mul_b2/fa1_c1_r[19] , \mul_b2/fa1_c1_r[18] ,
         \mul_b2/fa1_c1_r[17] , \mul_b2/fa1_c1_r[16] , \mul_b2/fa1_c1_r[15] ,
         \mul_b2/fa1_c1_r[14] , \mul_b2/fa1_c1_r[13] , \mul_b2/fa1_c1_r[12] ,
         \mul_b2/fa1_c1_r[11] , \mul_b2/fa1_c1_r[10] , \mul_b2/fa1_c1_r[9] ,
         \mul_b2/fa1_s1_r[33] , \mul_b2/fa1_s1_r[32] , \mul_b2/fa1_s1_r[31] ,
         \mul_b2/fa1_s1_r[30] , \mul_b2/fa1_s1_r[29] , \mul_b2/fa1_s1_r[28] ,
         \mul_b2/fa1_s1_r[27] , \mul_b2/fa1_s1_r[26] , \mul_b2/fa1_s1_r[25] ,
         \mul_b2/fa1_s1_r[24] , \mul_b2/fa1_s1_r[23] , \mul_b2/fa1_s1_r[22] ,
         \mul_b2/fa1_s1_r[21] , \mul_b2/fa1_s1_r[20] , \mul_b2/fa1_s1_r[19] ,
         \mul_b2/fa1_s1_r[18] , \mul_b2/fa1_s1_r[17] , \mul_b2/fa1_s1_r[16] ,
         \mul_b2/fa1_s1_r[15] , \mul_b2/fa1_s1_r[14] , \mul_b2/fa1_s1_r[13] ,
         \mul_b2/fa1_s1_r[12] , \mul_b2/fa1_s1_r[11] , \mul_b2/fa1_s1_r[10] ,
         \mul_b2/fa1_s1_r[9] , \mul_b2/fa1_s1_r[8] , \mul_b2/fa1_s1_r[7] ,
         \mul_b2/fa1_s1_r[6] , \mul_b2/fa1_c0_r[32] , \mul_b2/fa1_c0_r[31] ,
         \mul_b2/fa1_c0_r[30] , \mul_b2/fa1_c0_r[29] , \mul_b2/fa1_c0_r[28] ,
         \mul_b2/fa1_c0_r[27] , \mul_b2/fa1_c0_r[26] , \mul_b2/fa1_c0_r[25] ,
         \mul_b2/fa1_c0_r[24] , \mul_b2/fa1_c0_r[23] , \mul_b2/fa1_c0_r[22] ,
         \mul_b2/fa1_c0_r[21] , \mul_b2/fa1_c0_r[20] , \mul_b2/fa1_c0_r[19] ,
         \mul_b2/fa1_c0_r[18] , \mul_b2/fa1_c0_r[17] , \mul_b2/fa1_c0_r[16] ,
         \mul_b2/fa1_c0_r[15] , \mul_b2/fa1_c0_r[14] , \mul_b2/fa1_c0_r[13] ,
         \mul_b2/fa1_c0_r[12] , \mul_b2/fa1_c0_r[11] , \mul_b2/fa1_c0_r[10] ,
         \mul_b2/fa1_c0_r[9] , \mul_b2/fa1_c0_r[8] , \mul_b2/fa1_c0_r[7] ,
         \mul_b2/fa1_c0_r[6] , \mul_b2/fa1_c0_r[5] , \mul_b2/fa1_c0_r[4] ,
         \mul_b2/fa1_c0_r[3] , \mul_b2/fa1_s0_r[33] , \mul_b2/fa1_s0_r[32] ,
         \mul_b2/fa1_s0_r[31] , \mul_b2/fa1_s0_r[30] , \mul_b2/fa1_s0_r[29] ,
         \mul_b2/fa1_s0_r[28] , \mul_b2/fa1_s0_r[27] , \mul_b2/fa1_s0_r[26] ,
         \mul_b2/fa1_s0_r[25] , \mul_b2/fa1_s0_r[24] , \mul_b2/fa1_s0_r[23] ,
         \mul_b2/fa1_s0_r[22] , \mul_b2/fa1_s0_r[21] , \mul_b2/fa1_s0_r[20] ,
         \mul_b2/fa1_s0_r[19] , \mul_b2/fa1_s0_r[18] , \mul_b2/fa1_s0_r[17] ,
         \mul_b2/fa1_s0_r[16] , \mul_b2/fa1_s0_r[15] , \mul_b2/fa1_s0_r[14] ,
         \mul_b2/fa1_s0_r[13] , \mul_b2/fa1_s0_r[12] , \mul_b2/fa1_s0_r[11] ,
         \mul_b2/fa1_s0_r[10] , \mul_b2/fa1_s0_r[9] , \mul_b2/fa1_s0_r[8] ,
         \mul_b2/fa1_s0_r[7] , \mul_b2/fa1_s0_r[6] , \mul_b2/fa1_s0_r[5] ,
         \mul_b2/fa1_s0_r[4] , \mul_b2/fa1_c1[23] , \mul_b2/fa1_c1[22] ,
         \mul_b2/fa1_c1[21] , \mul_b2/fa1_c1[20] , \mul_b2/fa1_c1[19] ,
         \mul_b2/fa1_c1[18] , \mul_b2/fa1_c1[17] , \mul_b2/fa1_c1[16] ,
         \mul_b2/fa1_c1[15] , \mul_b2/fa1_c1[14] , \mul_b2/fa1_c1[13] ,
         \mul_b2/fa1_c1[12] , \mul_b2/fa1_c1[11] , \mul_b2/fa1_c1[10] ,
         \mul_b2/fa1_c1[9] , \mul_b2/fa1_s1[28] , \mul_b2/fa1_s1[23] ,
         \mul_b2/fa1_s1[22] , \mul_b2/fa1_s1[21] , \mul_b2/fa1_s1[20] ,
         \mul_b2/fa1_s1[19] , \mul_b2/fa1_s1[18] , \mul_b2/fa1_s1[17] ,
         \mul_b2/fa1_s1[16] , \mul_b2/fa1_s1[15] , \mul_b2/fa1_s1[14] ,
         \mul_b2/fa1_s1[13] , \mul_b2/fa1_s1[12] , \mul_b2/fa1_s1[11] ,
         \mul_b2/fa1_s1[10] , \mul_b2/fa1_s1[9] , \mul_b2/fa1_s1[7] ,
         \mul_b2/fa1_c0[18] , \mul_b2/fa1_c0[17] , \mul_b2/fa1_c0[16] ,
         \mul_b2/fa1_c0[15] , \mul_b2/fa1_c0[14] , \mul_b2/fa1_c0[13] ,
         \mul_b2/fa1_c0[12] , \mul_b2/fa1_c0[11] , \mul_b2/fa1_c0[10] ,
         \mul_b2/fa1_c0[9] , \mul_b2/fa1_c0[8] , \mul_b2/fa1_c0[7] ,
         \mul_b2/fa1_c0[6] , \mul_b2/fa1_c0[5] , \mul_b2/fa1_c0[4] ,
         \mul_b2/fa1_c0[3] , \mul_b2/fa1_s0[18] , \mul_b2/fa1_s0[17] ,
         \mul_b2/fa1_s0[16] , \mul_b2/fa1_s0[15] , \mul_b2/fa1_s0[14] ,
         \mul_b2/fa1_s0[13] , \mul_b2/fa1_s0[12] , \mul_b2/fa1_s0[11] ,
         \mul_b2/fa1_s0[10] , \mul_b2/fa1_s0[9] , \mul_b2/fa1_s0[8] ,
         \mul_b2/fa1_s0[7] , \mul_b2/fa1_s0[6] , \mul_b2/fa1_s0[5] ,
         \mul_b2/fa1_s0[4] , \mul_a1/result_sat[15] , \mul_a1/result_sat[14] ,
         \mul_a1/result_sat[13] , \mul_a1/result_sat[12] ,
         \mul_a1/result_sat[11] , \mul_a1/result_sat[10] ,
         \mul_a1/result_sat[9] , \mul_a1/result_sat[8] ,
         \mul_a1/result_sat[7] , \mul_a1/result_sat[6] ,
         \mul_a1/result_sat[5] , \mul_a1/result_sat[4] ,
         \mul_a1/result_sat[3] , \mul_a1/result_sat[2] ,
         \mul_a1/result_sat[1] , \mul_a1/result_sat[0] , \mul_a1/fa1_s2_r[33] ,
         \mul_a1/fa1_s2_r[32] , \mul_a1/fa1_s2_r[31] , \mul_a1/fa1_s2_r[30] ,
         \mul_a1/fa1_s2_r[29] , \mul_a1/fa1_s2_r[28] , \mul_a1/fa1_s2_r[27] ,
         \mul_a1/fa1_s2_r[26] , \mul_a1/fa1_s2_r[25] , \mul_a1/fa1_s2_r[24] ,
         \mul_a1/fa1_s2_r[23] , \mul_a1/fa1_s2_r[22] , \mul_a1/fa1_s2_r[21] ,
         \mul_a1/fa1_s2_r[20] , \mul_a1/fa1_s2_r[19] , \mul_a1/fa1_s2_r[18] ,
         \mul_a1/fa1_s2_r[17] , \mul_a1/fa1_s2_r[16] , \mul_a1/fa1_s2_r[15] ,
         \mul_a1/fa1_s2_r[14] , \mul_a1/fa1_c1_r[32] , \mul_a1/fa1_c1_r[31] ,
         \mul_a1/fa1_c1_r[30] , \mul_a1/fa1_c1_r[29] , \mul_a1/fa1_c1_r[28] ,
         \mul_a1/fa1_c1_r[27] , \mul_a1/fa1_c1_r[26] , \mul_a1/fa1_c1_r[25] ,
         \mul_a1/fa1_c1_r[24] , \mul_a1/fa1_c1_r[23] , \mul_a1/fa1_c1_r[22] ,
         \mul_a1/fa1_c1_r[21] , \mul_a1/fa1_c1_r[20] , \mul_a1/fa1_c1_r[19] ,
         \mul_a1/fa1_c1_r[18] , \mul_a1/fa1_c1_r[17] , \mul_a1/fa1_c1_r[16] ,
         \mul_a1/fa1_c1_r[15] , \mul_a1/fa1_c1_r[14] , \mul_a1/fa1_c1_r[13] ,
         \mul_a1/fa1_c1_r[12] , \mul_a1/fa1_c1_r[11] , \mul_a1/fa1_c1_r[10] ,
         \mul_a1/fa1_c1_r[9] , \mul_a1/fa1_c1_r[8] , \mul_a1/fa1_s1_r[33] ,
         \mul_a1/fa1_s1_r[32] , \mul_a1/fa1_s1_r[31] , \mul_a1/fa1_s1_r[30] ,
         \mul_a1/fa1_s1_r[29] , \mul_a1/fa1_s1_r[28] , \mul_a1/fa1_s1_r[27] ,
         \mul_a1/fa1_s1_r[26] , \mul_a1/fa1_s1_r[25] , \mul_a1/fa1_s1_r[24] ,
         \mul_a1/fa1_s1_r[23] , \mul_a1/fa1_s1_r[22] , \mul_a1/fa1_s1_r[21] ,
         \mul_a1/fa1_s1_r[20] , \mul_a1/fa1_s1_r[19] , \mul_a1/fa1_s1_r[18] ,
         \mul_a1/fa1_s1_r[17] , \mul_a1/fa1_s1_r[16] , \mul_a1/fa1_s1_r[15] ,
         \mul_a1/fa1_s1_r[14] , \mul_a1/fa1_s1_r[13] , \mul_a1/fa1_s1_r[12] ,
         \mul_a1/fa1_s1_r[11] , \mul_a1/fa1_s1_r[10] , \mul_a1/fa1_s1_r[9] ,
         \mul_a1/fa1_s1_r[8] , \mul_a1/fa1_s1_r[7] , \mul_a1/fa1_s0_r[33] ,
         \mul_a1/fa1_s0_r[32] , \mul_a1/fa1_s0_r[31] , \mul_a1/fa1_s0_r[30] ,
         \mul_a1/fa1_s0_r[29] , \mul_a1/fa1_s0_r[28] , \mul_a1/fa1_s0_r[27] ,
         \mul_a1/fa1_s0_r[26] , \mul_a1/fa1_s0_r[25] , \mul_a1/fa1_s0_r[24] ,
         \mul_a1/fa1_s0_r[23] , \mul_a1/fa1_s0_r[22] , \mul_a1/fa1_s0_r[21] ,
         \mul_a1/fa1_s0_r[20] , \mul_a1/fa1_s0_r[19] , \mul_a1/fa1_s0_r[18] ,
         \mul_a1/fa1_s0_r[17] , \mul_a1/fa1_s0_r[16] , \mul_a1/fa1_s0_r[15] ,
         \mul_a1/fa1_s0_r[14] , \mul_a1/fa1_s0_r[13] , \mul_a1/fa1_s0_r[12] ,
         \mul_a1/fa1_s0_r[11] , \mul_a1/fa1_s0_r[10] , \mul_a1/fa1_s0_r[9] ,
         \mul_a1/fa1_s0_r[8] , \mul_a1/fa1_s0_r[7] , \mul_a1/fa1_c1[22] ,
         \mul_a1/fa1_c1[21] , \mul_a1/fa1_c1[20] , \mul_a1/fa1_c1[19] ,
         \mul_a1/fa1_c1[18] , \mul_a1/fa1_c1[17] , \mul_a1/fa1_c1[16] ,
         \mul_a1/fa1_c1[15] , \mul_a1/fa1_c1[14] , \mul_a1/fa1_c1[13] ,
         \mul_a1/fa1_c1[12] , \mul_a1/fa1_c1[11] , \mul_a1/fa1_c1[10] ,
         \mul_a1/fa1_c1[9] , \mul_a1/fa1_c1[8] , \mul_a1/fa1_s1[22] ,
         \mul_a1/fa1_s1[21] , \mul_a1/fa1_s1[20] , \mul_a1/fa1_s1[19] ,
         \mul_a1/fa1_s1[18] , \mul_a1/fa1_s1[17] , \mul_a1/fa1_s1[16] ,
         \mul_a1/fa1_s1[15] , \mul_a1/fa1_s1[14] , \mul_a1/fa1_s1[13] ,
         \mul_a1/fa1_s1[12] , \mul_a1/fa1_s1[11] , \mul_a1/fa1_s1[10] ,
         \mul_a1/fa1_s1[9] , \mul_a1/fa1_s1[8] , \mul_a1/fa1_s1[7] ,
         \mul_a2/result_sat[15] , \mul_a2/result_sat[14] ,
         \mul_a2/result_sat[13] , \mul_a2/result_sat[12] ,
         \mul_a2/result_sat[11] , \mul_a2/result_sat[10] ,
         \mul_a2/result_sat[9] , \mul_a2/result_sat[8] ,
         \mul_a2/result_sat[7] , \mul_a2/result_sat[6] ,
         \mul_a2/result_sat[5] , \mul_a2/result_sat[4] ,
         \mul_a2/result_sat[3] , \mul_a2/result_sat[2] ,
         \mul_a2/result_sat[1] , \mul_a2/result_sat[0] , \mul_a2/fa1_s2_r[33] ,
         \mul_a2/fa1_s2_r[32] , \mul_a2/fa1_s2_r[31] , \mul_a2/fa1_s2_r[30] ,
         \mul_a2/fa1_s2_r[29] , \mul_a2/fa1_s2_r[28] , \mul_a2/fa1_s2_r[27] ,
         \mul_a2/fa1_s2_r[26] , \mul_a2/fa1_s2_r[25] , \mul_a2/fa1_s2_r[24] ,
         \mul_a2/fa1_s2_r[23] , \mul_a2/fa1_s2_r[22] , \mul_a2/fa1_s2_r[21] ,
         \mul_a2/fa1_s2_r[20] , \mul_a2/fa1_s2_r[19] , \mul_a2/fa1_s2_r[18] ,
         \mul_a2/fa1_s2_r[17] , \mul_a2/fa1_s2_r[16] , \mul_a2/fa1_s2_r[15] ,
         \mul_a2/fa1_s2_r[14] , \mul_a2/fa1_s2_r[13] , \mul_a2/fa1_s1_r[33] ,
         \mul_a2/fa1_s1_r[32] , \mul_a2/fa1_s1_r[31] , \mul_a2/fa1_s1_r[30] ,
         \mul_a2/fa1_s1_r[29] , \mul_a2/fa1_s1_r[28] , \mul_a2/fa1_s1_r[27] ,
         \mul_a2/fa1_s1_r[26] , \mul_a2/fa1_s1_r[25] , \mul_a2/fa1_s1_r[24] ,
         \mul_a2/fa1_s1_r[23] , \mul_a2/fa1_s1_r[22] , \mul_a2/fa1_s1_r[21] ,
         \mul_a2/fa1_s1_r[20] , \mul_a2/fa1_s1_r[19] , \mul_a2/fa1_s1_r[18] ,
         \mul_a2/fa1_s1_r[17] , \mul_a2/fa1_s1_r[16] , \mul_a2/fa1_s1_r[15] ,
         \mul_a2/fa1_s1_r[14] , \mul_a2/fa1_s1_r[13] , \mul_a2/fa1_s1_r[12] ,
         \mul_a2/fa1_s1_r[11] , \mul_a2/fa1_c0_r[16] , \mul_a2/fa1_c0_r[15] ,
         \mul_a2/fa1_c0_r[14] , \mul_a2/fa1_c0_r[13] , \mul_a2/fa1_c0_r[12] ,
         \mul_a2/fa1_c0_r[11] , \mul_a2/fa1_c0_r[10] , \mul_a2/fa1_c0_r[9] ,
         \mul_a2/fa1_c0_r[8] , \mul_a2/fa1_c0_r[7] , \mul_a2/fa1_c0_r[6] ,
         \mul_a2/fa1_c0_r[5] , \mul_a2/fa1_c0_r[4] , \mul_a2/fa1_c0_r[3] ,
         \mul_a2/fa1_c0_r[2] , \mul_a2/fa1_s0_r[33] , \mul_a2/fa1_s0_r[32] ,
         \mul_a2/fa1_s0_r[31] , \mul_a2/fa1_s0_r[30] , \mul_a2/fa1_s0_r[29] ,
         \mul_a2/fa1_s0_r[28] , \mul_a2/fa1_s0_r[27] , \mul_a2/fa1_s0_r[26] ,
         \mul_a2/fa1_s0_r[25] , \mul_a2/fa1_s0_r[24] , \mul_a2/fa1_s0_r[23] ,
         \mul_a2/fa1_s0_r[22] , \mul_a2/fa1_s0_r[21] , \mul_a2/fa1_s0_r[20] ,
         \mul_a2/fa1_s0_r[19] , \mul_a2/fa1_s0_r[18] , \mul_a2/fa1_s0_r[17] ,
         \mul_a2/fa1_s0_r[16] , \mul_a2/fa1_s0_r[15] , \mul_a2/fa1_s0_r[14] ,
         \mul_a2/fa1_s0_r[13] , \mul_a2/fa1_s0_r[12] , \mul_a2/fa1_s0_r[11] ,
         \mul_a2/fa1_s0_r[10] , \mul_a2/fa1_s0_r[9] , \mul_a2/fa1_s0_r[8] ,
         \mul_a2/fa1_s0_r[7] , \mul_a2/fa1_s0_r[6] , \mul_a2/fa1_s0_r[5] ,
         \mul_a2/fa1_s0_r[4] , \mul_a2/fa1_s0_r[3] , \mul_a2/fa1_c0[16] ,
         \mul_a2/fa1_c0[15] , \mul_a2/fa1_c0[14] , \mul_a2/fa1_c0[13] ,
         \mul_a2/fa1_c0[12] , \mul_a2/fa1_c0[11] , \mul_a2/fa1_c0[10] ,
         \mul_a2/fa1_c0[9] , \mul_a2/fa1_c0[8] , \mul_a2/fa1_c0[7] ,
         \mul_a2/fa1_c0[6] , \mul_a2/fa1_c0[5] , \mul_a2/fa1_c0[4] ,
         \mul_a2/fa1_c0[3] , \mul_a2/fa1_c0[2] , \mul_a2/fa1_s0[31] ,
         \mul_a2/fa1_s0[16] , \mul_a2/fa1_s0[15] , \mul_a2/fa1_s0[14] ,
         \mul_a2/fa1_s0[13] , \mul_a2/fa1_s0[12] , \mul_a2/fa1_s0[11] ,
         \mul_a2/fa1_s0[10] , \mul_a2/fa1_s0[9] , \mul_a2/fa1_s0[8] ,
         \mul_a2/fa1_s0[7] , \mul_a2/fa1_s0[6] , \mul_a2/fa1_s0[5] ,
         \mul_a2/fa1_s0[4] , \mul_a2/fa1_s0[3] , \C63/DATA4_12 ,
         \C63/DATA4_13 , \C63/DATA4_14 , \C63/DATA4_15 , \C63/DATA4_16 ,
         \C63/DATA4_17 , \C63/DATA4_18 , \C63/DATA4_19 , \C63/DATA4_20 ,
         \C63/DATA4_21 , \C63/DATA4_22 , \C63/DATA4_23 , \C63/DATA4_24 ,
         \C63/DATA4_25 , \C63/DATA4_26 , \C56/DATA4_15 , \C56/DATA4_16 ,
         \C56/DATA4_17 , \C56/DATA4_18 , \C56/DATA4_19 , \C56/DATA4_20 ,
         \C56/DATA4_21 , \C56/DATA4_22 , \C56/DATA4_23 , \C56/DATA4_24 ,
         \C56/DATA4_25 , \C56/DATA4_26 , \C56/DATA4_27 , \C56/DATA4_28 ,
         \C56/DATA4_29 , \C56/DATA4_30 , \C49/DATA3_7 , \C49/DATA3_8 ,
         \C49/DATA3_9 , \C49/DATA3_10 , \C49/DATA3_11 , \C49/DATA3_12 ,
         \C49/DATA3_13 , \C49/DATA3_14 , \C49/DATA3_15 , \C49/DATA3_16 ,
         \C43/DATA4_8 , \C33/DATA4_17 , \C33/DATA4_18 , \C33/DATA4_19 ,
         \C33/DATA4_20 , \DP_OP_331J1_157_5454/n87 ,
         \DP_OP_371J1_181_1383/n79 , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917;
  wire   [15:0] x_z1;
  wire   [15:0] x_z2;
  wire   [15:0] y_z1;
  wire   [15:0] y_z2;
  wire   [15:0] x_reg2;
  wire   [15:0] p_b0;
  wire   [15:0] p_b1;
  wire   [15:0] p_b2;
  wire   [15:0] p_a1;
  wire   [15:0] p_a2;

  HS65_GS_DFPRQX4 valid_T1_reg ( .D(n1821), .CP(clk), .RN(rst_n), .Q(valid_T1)
         );
  HS65_GS_DFPRQX4 valid_T2_reg ( .D(valid_T1), .CP(clk), .RN(rst_n), .Q(
        valid_T2) );
  HS65_GS_DFPRQX4 valid_T3_reg ( .D(valid_T2), .CP(clk), .RN(rst_n), .Q(
        valid_T3) );
  HS65_GS_DFPRQX4 valid_out_reg ( .D(valid_T3), .CP(clk), .RN(rst_n), .Q(
        valid_out) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[0]  ( .D(\mul_b0/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[0]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[1]  ( .D(\mul_b0/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[1]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[2]  ( .D(\mul_b0/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[2]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[3]  ( .D(\mul_b0/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[3]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[4]  ( .D(\mul_b0/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[4]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[5]  ( .D(\mul_b0/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[5]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[6]  ( .D(\mul_b0/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[6]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[7]  ( .D(\mul_b0/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[7]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[8]  ( .D(\mul_b0/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[8]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[9]  ( .D(\mul_b0/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[9]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[10]  ( .D(\mul_b0/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[10]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[11]  ( .D(\mul_b0/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[11]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[12]  ( .D(\mul_b0/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[12]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[13]  ( .D(\mul_b0/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[13]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[14]  ( .D(\mul_b0/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[14]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[15]  ( .D(\mul_b0/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[15]) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[12]  ( .D(x_z1[0]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[13]  ( .D(x_z1[1]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[14]  ( .D(x_z1[2]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[15]  ( .D(x_z1[3]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[16]  ( .D(x_z1[4]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[17]  ( .D(x_z1[5]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[18]  ( .D(x_z1[6]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[19]  ( .D(x_z1[7]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[20]  ( .D(x_z1[8]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[21]  ( .D(x_z1[9]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[22]  ( .D(x_z1[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[23]  ( .D(x_z1[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[24]  ( .D(x_z1[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[25]  ( .D(x_z1[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[26]  ( .D(x_z1[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[27]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[28]  ( .D(n1820), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[29]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[30]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[31]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[32]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[33]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[8]  ( .D(x_z1[0]), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[9]  ( .D(x_z1[1]), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[10]  ( .D(x_z1[2]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[11]  ( .D(x_z1[3]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[12]  ( .D(x_z1[4]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[13]  ( .D(x_z1[5]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[14]  ( .D(x_z1[6]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[15]  ( .D(x_z1[7]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[16]  ( .D(x_z1[8]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[17]  ( .D(x_z1[9]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[18]  ( .D(x_z1[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[19]  ( .D(x_z1[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[20]  ( .D(x_z1[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[21]  ( .D(x_z1[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[22]  ( .D(x_z1[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[23]  ( .D(n1820), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[24]  ( .D(n1820), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[25]  ( .D(n1820), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[26]  ( .D(n1820), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[27]  ( .D(n1820), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[28]  ( .D(n1820), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[29]  ( .D(n1820), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[30]  ( .D(n1820), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[31]  ( .D(n1820), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[32]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[33]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[5]  ( .D(\mul_b0/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[6]  ( .D(\mul_b0/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[7]  ( .D(\mul_b0/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[8]  ( .D(\mul_b0/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[9]  ( .D(\mul_b0/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[10]  ( .D(\mul_b0/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[11]  ( .D(\mul_b0/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[12]  ( .D(\mul_b0/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[13]  ( .D(\mul_b0/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[14]  ( .D(\mul_b0/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[15]  ( .D(\mul_b0/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[16]  ( .D(\mul_b0/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[17]  ( .D(\mul_b0/fa1_c0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[18]  ( .D(\mul_b0/fa1_c0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[19]  ( .D(\mul_b0/fa1_c0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[20]  ( .D(\mul_b0/fa1_c0[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[6]  ( .D(\mul_b0/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[7]  ( .D(\mul_b0/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[8]  ( .D(\mul_b0/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[9]  ( .D(\mul_b0/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[10]  ( .D(\mul_b0/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[11]  ( .D(\mul_b0/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[12]  ( .D(\mul_b0/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[13]  ( .D(\mul_b0/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[14]  ( .D(\mul_b0/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[15]  ( .D(\mul_b0/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[16]  ( .D(\mul_b0/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[17]  ( .D(\mul_b0/fa1_s0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[18]  ( .D(\mul_b0/fa1_s0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[19]  ( .D(\mul_b0/fa1_s0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[20]  ( .D(\mul_b0/fa1_s0[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[21]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[22]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[23]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[24]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[25]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[26]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[27]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[28]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[29]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[30]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[31]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[32]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[33]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[0]  ( .D(\mul_b1/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[0]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[1]  ( .D(\mul_b1/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[1]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[2]  ( .D(\mul_b1/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[2]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[3]  ( .D(\mul_b1/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[3]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[4]  ( .D(\mul_b1/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[4]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[5]  ( .D(\mul_b1/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[5]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[6]  ( .D(\mul_b1/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[6]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[7]  ( .D(\mul_b1/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[7]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[8]  ( .D(\mul_b1/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[8]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[9]  ( .D(\mul_b1/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[9]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[10]  ( .D(\mul_b1/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[10]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[11]  ( .D(\mul_b1/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[11]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[12]  ( .D(\mul_b1/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[12]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[13]  ( .D(\mul_b1/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[13]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[14]  ( .D(\mul_b1/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[14]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[15]  ( .D(\mul_b1/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[15]) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[13]  ( .D(x_z2[0]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[14]  ( .D(\mul_b1/fa1_s2[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[15]  ( .D(\mul_b1/fa1_s2[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[16]  ( .D(\mul_b1/fa1_s2[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[17]  ( .D(\mul_b1/fa1_s2[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[18]  ( .D(\mul_b1/fa1_s2[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[19]  ( .D(\mul_b1/fa1_s2[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[20]  ( .D(\mul_b1/fa1_s2[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[21]  ( .D(\mul_b1/fa1_s2[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[22]  ( .D(\mul_b1/fa1_s2[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[23]  ( .D(\mul_b1/fa1_s2[23] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[24]  ( .D(\mul_b1/fa1_s2[24] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[25]  ( .D(\mul_b1/fa1_s2[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[26]  ( .D(\mul_b1/fa1_s2[26] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[27]  ( .D(\mul_b1/fa1_s2[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[28]  ( .D(\mul_b1/fa1_s2[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[29]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[30]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[31]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[32]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[33]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[8]  ( .D(\mul_b1/fa1_c1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[9]  ( .D(\mul_b1/fa1_c1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[10]  ( .D(\mul_b1/fa1_c1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[11]  ( .D(\mul_b1/fa1_c1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[12]  ( .D(\mul_b1/fa1_c1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[13]  ( .D(\mul_b1/fa1_c1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[14]  ( .D(\mul_b1/fa1_c1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[15]  ( .D(\mul_b1/fa1_c1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[16]  ( .D(\mul_b1/fa1_c1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[17]  ( .D(\mul_b1/fa1_c1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[18]  ( .D(\mul_b1/fa1_c1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[19]  ( .D(\mul_b1/fa1_c1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[20]  ( .D(\mul_b1/fa1_c1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[21]  ( .D(\mul_b1/fa1_c1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[22]  ( .D(\mul_b1/fa1_c1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[23]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[24]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[25]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[26]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[27]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[28]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[29]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[30]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[31]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[32]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[6]  ( .D(x_z2[0]), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s1_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[7]  ( .D(\mul_b1/fa1_s1[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s1_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[8]  ( .D(\mul_b1/fa1_s1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[9]  ( .D(\mul_b1/fa1_s1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[10]  ( .D(\mul_b1/fa1_s1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[11]  ( .D(\mul_b1/fa1_s1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[12]  ( .D(\mul_b1/fa1_s1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[13]  ( .D(\mul_b1/fa1_s1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[14]  ( .D(\mul_b1/fa1_s1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[15]  ( .D(\mul_b1/fa1_s1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[16]  ( .D(\mul_b1/fa1_s1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[17]  ( .D(\mul_b1/fa1_s1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[18]  ( .D(\mul_b1/fa1_s1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[19]  ( .D(\mul_b1/fa1_s1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[20]  ( .D(\mul_b1/fa1_s1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[21]  ( .D(\mul_b1/fa1_s1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[22]  ( .D(\mul_b1/fa1_s1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[23]  ( .D(\mul_b1/fa1_s1[23] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[24]  ( .D(\mul_b1/fa1_s1[24] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[25]  ( .D(\mul_b1/fa1_s1[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[26]  ( .D(\mul_b1/fa1_s1[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[27]  ( .D(\mul_b1/fa1_s1[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[28]  ( .D(\mul_b1/fa1_s1[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[29]  ( .D(\mul_b1/fa1_s1[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[30]  ( .D(\mul_b1/fa1_s1[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[31]  ( .D(\mul_b1/fa1_s1[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[32]  ( .D(\mul_b1/fa1_s1[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[33]  ( .D(\mul_b1/fa1_s1[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[2]  ( .D(n1816), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[2] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[3]  ( .D(n1818), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[3] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[4]  ( .D(n1817), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[5]  ( .D(\mul_b1/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[6]  ( .D(\mul_b1/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[7]  ( .D(\mul_b1/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[8]  ( .D(\mul_b1/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[9]  ( .D(\mul_b1/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[10]  ( .D(\mul_b1/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[11]  ( .D(\mul_b1/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[12]  ( .D(\mul_b1/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[13]  ( .D(\mul_b1/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[14]  ( .D(\mul_b1/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[15]  ( .D(\mul_b1/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[16]  ( .D(\mul_b1/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[17]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_c0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[18]  ( .D(\DP_OP_331J1_157_5454/n87 ), 
        .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[19]  ( .D(\DP_OP_331J1_157_5454/n87 ), 
        .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[20]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_c0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[21]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_c0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[22]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_c0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[23]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_c0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[24]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_c0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[25]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_c0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[26]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_c0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[27]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_c0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[28]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_c0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[29]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_c0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[30]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_c0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[31]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_c0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[32]  ( .D(\DP_OP_331J1_157_5454/n87 ), 
        .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[3]  ( .D(\mul_b1/fa1_s0[3] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[3] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[4]  ( .D(\mul_b1/fa1_s0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[5]  ( .D(\mul_b1/fa1_s0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[6]  ( .D(\mul_b1/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[7]  ( .D(\mul_b1/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[8]  ( .D(\mul_b1/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[9]  ( .D(\mul_b1/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[10]  ( .D(\mul_b1/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[11]  ( .D(\mul_b1/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[12]  ( .D(\mul_b1/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[13]  ( .D(\mul_b1/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[14]  ( .D(\mul_b1/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[15]  ( .D(\mul_b1/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[16]  ( .D(\mul_b1/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[17]  ( .D(\C33/DATA4_17 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[18]  ( .D(\C33/DATA4_18 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[19]  ( .D(\C33/DATA4_19 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[20]  ( .D(\C33/DATA4_20 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[21]  ( .D(n1813), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[22]  ( .D(n1813), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[23]  ( .D(n1813), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[24]  ( .D(n1813), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[25]  ( .D(n1813), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[26]  ( .D(n1813), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[27]  ( .D(n1813), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[28]  ( .D(n1813), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[29]  ( .D(n1813), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[30]  ( .D(n1813), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[31]  ( .D(n1813), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[32]  ( .D(n1813), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[33]  ( .D(n1813), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[14]  ( .D(\mul_b1/fa1_c2[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[15]  ( .D(\mul_b1/fa1_c2[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[16]  ( .D(\mul_b1/fa1_c2[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[17]  ( .D(\mul_b1/fa1_c2[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[18]  ( .D(\mul_b1/fa1_c2[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[19]  ( .D(\mul_b1/fa1_c2[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[20]  ( .D(\mul_b1/fa1_c2[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[21]  ( .D(\mul_b1/fa1_c2[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[22]  ( .D(\mul_b1/fa1_c2[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[23]  ( .D(\mul_b1/fa1_c2[23] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[24]  ( .D(\mul_b1/fa1_c2[24] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[25]  ( .D(\mul_b1/fa1_c2[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[26]  ( .D(\mul_b1/fa1_c2[26] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[27]  ( .D(\mul_b1/fa1_c2[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[28]  ( .D(\mul_b1/fa1_c2[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[0]  ( .D(\mul_b2/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[0]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[1]  ( .D(\mul_b2/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[1]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[2]  ( .D(\mul_b2/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[2]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[3]  ( .D(\mul_b2/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[3]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[4]  ( .D(\mul_b2/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[4]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[5]  ( .D(\mul_b2/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[5]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[6]  ( .D(\mul_b2/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[6]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[7]  ( .D(\mul_b2/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[7]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[8]  ( .D(\mul_b2/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[8]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[9]  ( .D(\mul_b2/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[9]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[10]  ( .D(\mul_b2/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[10]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[11]  ( .D(\mul_b2/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[11]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[12]  ( .D(\mul_b2/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[12]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[13]  ( .D(\mul_b2/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[13]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[14]  ( .D(\mul_b2/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[14]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[15]  ( .D(\mul_b2/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[15]) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[12]  ( .D(x_reg2[0]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[13]  ( .D(x_reg2[1]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[14]  ( .D(x_reg2[2]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[15]  ( .D(x_reg2[3]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[16]  ( .D(x_reg2[4]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[17]  ( .D(x_reg2[5]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[18]  ( .D(x_reg2[6]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[19]  ( .D(x_reg2[7]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[20]  ( .D(x_reg2[8]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[21]  ( .D(x_reg2[9]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[22]  ( .D(x_reg2[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[23]  ( .D(x_reg2[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[24]  ( .D(x_reg2[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[25]  ( .D(x_reg2[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[26]  ( .D(x_reg2[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[27]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[28]  ( .D(\DP_OP_371J1_181_1383/n79 ), 
        .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[29]  ( .D(\DP_OP_371J1_181_1383/n79 ), 
        .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[30]  ( .D(\DP_OP_371J1_181_1383/n79 ), 
        .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[31]  ( .D(\DP_OP_371J1_181_1383/n79 ), 
        .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[32]  ( .D(\DP_OP_371J1_181_1383/n79 ), 
        .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[33]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c1_r_reg[9]  ( .D(\mul_b2/fa1_c1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c1_r_reg[10]  ( .D(\mul_b2/fa1_c1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c1_r_reg[11]  ( .D(\mul_b2/fa1_c1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c1_r_reg[12]  ( .D(\mul_b2/fa1_c1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c1_r_reg[13]  ( .D(\mul_b2/fa1_c1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c1_r_reg[14]  ( .D(\mul_b2/fa1_c1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c1_r_reg[15]  ( .D(\mul_b2/fa1_c1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c1_r_reg[16]  ( .D(\mul_b2/fa1_c1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c1_r_reg[17]  ( .D(\mul_b2/fa1_c1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c1_r_reg[18]  ( .D(\mul_b2/fa1_c1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c1_r_reg[19]  ( .D(\mul_b2/fa1_c1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c1_r_reg[20]  ( .D(\mul_b2/fa1_c1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c1_r_reg[21]  ( .D(\mul_b2/fa1_c1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c1_r_reg[22]  ( .D(\mul_b2/fa1_c1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c1_r_reg[23]  ( .D(\mul_b2/fa1_c1[23] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[6]  ( .D(x_reg2[0]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[7]  ( .D(\mul_b2/fa1_s1[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[8]  ( .D(\C43/DATA4_8 ), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[9]  ( .D(\mul_b2/fa1_s1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[10]  ( .D(\mul_b2/fa1_s1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[11]  ( .D(\mul_b2/fa1_s1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[12]  ( .D(\mul_b2/fa1_s1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[13]  ( .D(\mul_b2/fa1_s1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[14]  ( .D(\mul_b2/fa1_s1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[15]  ( .D(\mul_b2/fa1_s1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[16]  ( .D(\mul_b2/fa1_s1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[17]  ( .D(\mul_b2/fa1_s1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[18]  ( .D(\mul_b2/fa1_s1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[19]  ( .D(\mul_b2/fa1_s1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[20]  ( .D(\mul_b2/fa1_s1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[21]  ( .D(\mul_b2/fa1_s1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[22]  ( .D(\mul_b2/fa1_s1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[23]  ( .D(\mul_b2/fa1_s1[23] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[24]  ( .D(\mul_b2/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[25]  ( .D(\mul_b2/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[26]  ( .D(\mul_b2/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[27]  ( .D(\mul_b2/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[28]  ( .D(\mul_b2/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[29]  ( .D(\mul_b2/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[30]  ( .D(\mul_b2/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[31]  ( .D(\mul_b2/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[32]  ( .D(\mul_b2/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[33]  ( .D(\mul_b2/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[3]  ( .D(\mul_b2/fa1_c0[3] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[3] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[4]  ( .D(\mul_b2/fa1_c0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[5]  ( .D(\mul_b2/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[6]  ( .D(\mul_b2/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[7]  ( .D(\mul_b2/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[8]  ( .D(\mul_b2/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[9]  ( .D(\mul_b2/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[10]  ( .D(\mul_b2/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[11]  ( .D(\mul_b2/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[12]  ( .D(\mul_b2/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[13]  ( .D(\mul_b2/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[14]  ( .D(\mul_b2/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[15]  ( .D(\mul_b2/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[16]  ( .D(\mul_b2/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[17]  ( .D(\mul_b2/fa1_c0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[18]  ( .D(\mul_b2/fa1_c0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[19]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[20]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[21]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[22]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[23]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[24]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[25]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[26]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[27]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[28]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[29]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[30]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[31]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[32]  ( .D(\DP_OP_371J1_181_1383/n79 ), 
        .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[4]  ( .D(\mul_b2/fa1_s0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[5]  ( .D(\mul_b2/fa1_s0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[6]  ( .D(\mul_b2/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[7]  ( .D(\mul_b2/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[8]  ( .D(\mul_b2/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[9]  ( .D(\mul_b2/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[10]  ( .D(\mul_b2/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[11]  ( .D(\mul_b2/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[12]  ( .D(\mul_b2/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[13]  ( .D(\mul_b2/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[14]  ( .D(\mul_b2/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[15]  ( .D(\mul_b2/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[16]  ( .D(\mul_b2/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[17]  ( .D(\mul_b2/fa1_s0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[18]  ( .D(\mul_b2/fa1_s0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[19]  ( .D(n1812), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[20]  ( .D(n1812), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[21]  ( .D(n1812), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[22]  ( .D(n1812), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[23]  ( .D(n1812), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[24]  ( .D(n1812), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[25]  ( .D(n1812), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[26]  ( .D(n1812), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[27]  ( .D(n1812), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[28]  ( .D(n1812), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[29]  ( .D(n1812), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[30]  ( .D(n1812), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[31]  ( .D(n1812), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[32]  ( .D(n1812), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[33]  ( .D(n1812), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[0]  ( .D(\mul_a1/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[0]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[1]  ( .D(\mul_a1/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[1]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[2]  ( .D(\mul_a1/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[2]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[3]  ( .D(\mul_a1/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[3]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[4]  ( .D(\mul_a1/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[4]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[5]  ( .D(\mul_a1/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[5]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[6]  ( .D(\mul_a1/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[6]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[7]  ( .D(\mul_a1/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[7]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[8]  ( .D(\mul_a1/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[8]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[9]  ( .D(\mul_a1/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[9]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[10]  ( .D(\mul_a1/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[10]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[11]  ( .D(\mul_a1/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[11]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[12]  ( .D(\mul_a1/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[12]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[13]  ( .D(\mul_a1/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[13]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[14]  ( .D(\mul_a1/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[14]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[15]  ( .D(\mul_a1/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[15]) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[14]  ( .D(\mul_a1/fa1_s1[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[15]  ( .D(\C56/DATA4_15 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[16]  ( .D(\C56/DATA4_16 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[17]  ( .D(\C56/DATA4_17 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[18]  ( .D(\C56/DATA4_18 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[19]  ( .D(\C56/DATA4_19 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[20]  ( .D(\C56/DATA4_20 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[21]  ( .D(\C56/DATA4_21 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[22]  ( .D(\C56/DATA4_22 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[23]  ( .D(\C56/DATA4_23 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[24]  ( .D(\C56/DATA4_24 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[25]  ( .D(\C56/DATA4_25 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[26]  ( .D(\C56/DATA4_26 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[27]  ( .D(\C56/DATA4_27 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[28]  ( .D(\C56/DATA4_28 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[29]  ( .D(\C56/DATA4_29 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[30]  ( .D(\C56/DATA4_30 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[31]  ( .D(n1815), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[32]  ( .D(n1815), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[33]  ( .D(n1815), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[8]  ( .D(\mul_a1/fa1_c1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_c1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[9]  ( .D(\mul_a1/fa1_c1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_c1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[10]  ( .D(\mul_a1/fa1_c1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[11]  ( .D(\mul_a1/fa1_c1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[12]  ( .D(\mul_a1/fa1_c1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[13]  ( .D(\mul_a1/fa1_c1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[14]  ( .D(\mul_a1/fa1_c1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[15]  ( .D(\mul_a1/fa1_c1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[16]  ( .D(\mul_a1/fa1_c1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[17]  ( .D(\mul_a1/fa1_c1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[18]  ( .D(\mul_a1/fa1_c1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[19]  ( .D(\mul_a1/fa1_c1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[20]  ( .D(\mul_a1/fa1_c1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[21]  ( .D(\mul_a1/fa1_c1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[22]  ( .D(\mul_a1/fa1_c1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[23]  ( .D(n1819), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_c1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[24]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_c1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[25]  ( .D(n1819), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_c1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[26]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_c1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[27]  ( .D(n1819), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_c1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[28]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_c1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[29]  ( .D(n1819), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_c1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[30]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_c1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[31]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_c1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[32]  ( .D(n1819), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_c1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[7]  ( .D(\mul_a1/fa1_s1[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[8]  ( .D(\mul_a1/fa1_s1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[9]  ( .D(\mul_a1/fa1_s1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[10]  ( .D(\mul_a1/fa1_s1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[11]  ( .D(\mul_a1/fa1_s1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[12]  ( .D(\mul_a1/fa1_s1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[13]  ( .D(\mul_a1/fa1_s1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[14]  ( .D(\mul_a1/fa1_s1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[15]  ( .D(\mul_a1/fa1_s1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[16]  ( .D(\mul_a1/fa1_s1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[17]  ( .D(\mul_a1/fa1_s1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[18]  ( .D(\mul_a1/fa1_s1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[19]  ( .D(\mul_a1/fa1_s1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[20]  ( .D(\mul_a1/fa1_s1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[21]  ( .D(\mul_a1/fa1_s1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[22]  ( .D(\mul_a1/fa1_s1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[23]  ( .D(y_z1[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[24]  ( .D(y_z1[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[25]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[26]  ( .D(n1819), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[27]  ( .D(n1819), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[28]  ( .D(n1819), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[29]  ( .D(n1819), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[30]  ( .D(n1819), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[31]  ( .D(n1819), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[32]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[33]  ( .D(n1819), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[7]  ( .D(\C49/DATA3_7 ), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[8]  ( .D(\C49/DATA3_8 ), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[9]  ( .D(\C49/DATA3_9 ), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[10]  ( .D(\C49/DATA3_10 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[11]  ( .D(\C49/DATA3_11 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[12]  ( .D(\C49/DATA3_12 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[13]  ( .D(\C49/DATA3_13 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[14]  ( .D(\C49/DATA3_14 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[15]  ( .D(\C49/DATA3_15 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[16]  ( .D(\C49/DATA3_16 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[17]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[18]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[19]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[20]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[21]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[22]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[23]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[24]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[25]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[26]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[27]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[28]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[29]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[30]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[31]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[32]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[33]  ( .D(n1811), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[0]  ( .D(\mul_a2/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[0]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[1]  ( .D(\mul_a2/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[1]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[2]  ( .D(\mul_a2/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[2]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[3]  ( .D(\mul_a2/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[3]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[4]  ( .D(\mul_a2/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[4]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[5]  ( .D(\mul_a2/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[5]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[6]  ( .D(\mul_a2/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[6]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[7]  ( .D(\mul_a2/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[7]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[8]  ( .D(\mul_a2/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[8]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[9]  ( .D(\mul_a2/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[9]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[10]  ( .D(\mul_a2/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[10]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[11]  ( .D(\mul_a2/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[11]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[12]  ( .D(\mul_a2/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[12]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[13]  ( .D(\mul_a2/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[13]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[14]  ( .D(\mul_a2/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[14]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[15]  ( .D(\mul_a2/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[15]) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[13]  ( .D(y_z2[0]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[14]  ( .D(y_z2[1]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[15]  ( .D(y_z2[2]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[16]  ( .D(y_z2[3]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[17]  ( .D(y_z2[4]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[18]  ( .D(y_z2[5]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[19]  ( .D(y_z2[6]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[20]  ( .D(y_z2[7]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[21]  ( .D(y_z2[8]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[22]  ( .D(y_z2[9]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[23]  ( .D(y_z2[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[24]  ( .D(y_z2[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[25]  ( .D(y_z2[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[26]  ( .D(y_z2[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[27]  ( .D(y_z2[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[28]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[29]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[30]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[31]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[32]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[33]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[11]  ( .D(y_z2[0]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[12]  ( .D(\C63/DATA4_12 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[13]  ( .D(\C63/DATA4_13 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[14]  ( .D(\C63/DATA4_14 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[15]  ( .D(\C63/DATA4_15 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[16]  ( .D(\C63/DATA4_16 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[17]  ( .D(\C63/DATA4_17 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[18]  ( .D(\C63/DATA4_18 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[19]  ( .D(\C63/DATA4_19 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[20]  ( .D(\C63/DATA4_20 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[21]  ( .D(\C63/DATA4_21 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[22]  ( .D(\C63/DATA4_22 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[23]  ( .D(\C63/DATA4_23 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[24]  ( .D(\C63/DATA4_24 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[25]  ( .D(\C63/DATA4_25 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[26]  ( .D(\C63/DATA4_26 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[27]  ( .D(n1814), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[28]  ( .D(n1814), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[29]  ( .D(n1814), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[30]  ( .D(n1814), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[31]  ( .D(n1814), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[32]  ( .D(n1814), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[33]  ( .D(n1814), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[2]  ( .D(\mul_a2/fa1_c0[2] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[2] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[3]  ( .D(\mul_a2/fa1_c0[3] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[3] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[4]  ( .D(\mul_a2/fa1_c0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[5]  ( .D(\mul_a2/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[6]  ( .D(\mul_a2/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[7]  ( .D(\mul_a2/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[8]  ( .D(\mul_a2/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[9]  ( .D(\mul_a2/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[10]  ( .D(\mul_a2/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[11]  ( .D(\mul_a2/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[12]  ( .D(\mul_a2/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[13]  ( .D(\mul_a2/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[14]  ( .D(\mul_a2/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[15]  ( .D(\mul_a2/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[16]  ( .D(\mul_a2/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[3]  ( .D(\mul_a2/fa1_s0[3] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[3] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[4]  ( .D(\mul_a2/fa1_s0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[5]  ( .D(\mul_a2/fa1_s0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[6]  ( .D(\mul_a2/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[7]  ( .D(\mul_a2/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[8]  ( .D(\mul_a2/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[9]  ( .D(\mul_a2/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[10]  ( .D(\mul_a2/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[11]  ( .D(\mul_a2/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[12]  ( .D(\mul_a2/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[13]  ( .D(\mul_a2/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[14]  ( .D(\mul_a2/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[15]  ( .D(\mul_a2/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[16]  ( .D(\mul_a2/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[17]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[18]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[19]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[20]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[21]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[22]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[23]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[24]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[25]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[26]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[27]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[28]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[29]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[30]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[31]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[32]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[33]  ( .D(\mul_a2/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \x_z1_reg[15]  ( .D(n1822), .CP(clk), .RN(rst_n), .Q(
        x_z1[15]) );
  HS65_GS_DFPRQX4 \x_z1_reg[14]  ( .D(n1823), .CP(clk), .RN(rst_n), .Q(
        x_z1[14]) );
  HS65_GS_DFPRQX4 \x_z1_reg[13]  ( .D(n1824), .CP(clk), .RN(rst_n), .Q(
        x_z1[13]) );
  HS65_GS_DFPRQX4 \x_z1_reg[12]  ( .D(n1825), .CP(clk), .RN(rst_n), .Q(
        x_z1[12]) );
  HS65_GS_DFPRQX4 \x_z1_reg[11]  ( .D(n1826), .CP(clk), .RN(rst_n), .Q(
        x_z1[11]) );
  HS65_GS_DFPRQX4 \x_z1_reg[10]  ( .D(n1827), .CP(clk), .RN(rst_n), .Q(
        x_z1[10]) );
  HS65_GS_DFPRQX4 \x_z1_reg[9]  ( .D(n1828), .CP(clk), .RN(rst_n), .Q(x_z1[9])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[8]  ( .D(n1829), .CP(clk), .RN(rst_n), .Q(x_z1[8])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[7]  ( .D(n1830), .CP(clk), .RN(rst_n), .Q(x_z1[7])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[6]  ( .D(n1831), .CP(clk), .RN(rst_n), .Q(x_z1[6])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[5]  ( .D(n1832), .CP(clk), .RN(rst_n), .Q(x_z1[5])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[4]  ( .D(n1833), .CP(clk), .RN(rst_n), .Q(x_z1[4])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[3]  ( .D(n1834), .CP(clk), .RN(rst_n), .Q(x_z1[3])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[2]  ( .D(n1835), .CP(clk), .RN(rst_n), .Q(x_z1[2])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[1]  ( .D(n1836), .CP(clk), .RN(rst_n), .Q(x_z1[1])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[0]  ( .D(n1837), .CP(clk), .RN(rst_n), .Q(x_z1[0])
         );
  HS65_GS_DFPRQX4 \x_z2_reg[15]  ( .D(n1838), .CP(clk), .RN(rst_n), .Q(
        x_z2[15]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[15]  ( .D(n1839), .CP(clk), .RN(rst_n), .Q(
        x_reg2[15]) );
  HS65_GS_DFPRQX4 \x_z2_reg[14]  ( .D(n1840), .CP(clk), .RN(rst_n), .Q(
        x_z2[14]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[14]  ( .D(n1841), .CP(clk), .RN(rst_n), .Q(
        x_reg2[14]) );
  HS65_GS_DFPRQX4 \x_z2_reg[13]  ( .D(n1842), .CP(clk), .RN(rst_n), .Q(
        x_z2[13]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[13]  ( .D(n1843), .CP(clk), .RN(rst_n), .Q(
        x_reg2[13]) );
  HS65_GS_DFPRQX4 \x_z2_reg[12]  ( .D(n1844), .CP(clk), .RN(rst_n), .Q(
        x_z2[12]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[12]  ( .D(n1845), .CP(clk), .RN(rst_n), .Q(
        x_reg2[12]) );
  HS65_GS_DFPRQX4 \x_z2_reg[11]  ( .D(n1846), .CP(clk), .RN(rst_n), .Q(
        x_z2[11]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[11]  ( .D(n1847), .CP(clk), .RN(rst_n), .Q(
        x_reg2[11]) );
  HS65_GS_DFPRQX4 \x_z2_reg[10]  ( .D(n1848), .CP(clk), .RN(rst_n), .Q(
        x_z2[10]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[10]  ( .D(n1849), .CP(clk), .RN(rst_n), .Q(
        x_reg2[10]) );
  HS65_GS_DFPRQX4 \x_z2_reg[9]  ( .D(n1850), .CP(clk), .RN(rst_n), .Q(x_z2[9])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[9]  ( .D(n1851), .CP(clk), .RN(rst_n), .Q(
        x_reg2[9]) );
  HS65_GS_DFPRQX4 \x_z2_reg[8]  ( .D(n1852), .CP(clk), .RN(rst_n), .Q(x_z2[8])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[8]  ( .D(n1853), .CP(clk), .RN(rst_n), .Q(
        x_reg2[8]) );
  HS65_GS_DFPRQX4 \x_z2_reg[7]  ( .D(n1854), .CP(clk), .RN(rst_n), .Q(x_z2[7])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[7]  ( .D(n1855), .CP(clk), .RN(rst_n), .Q(
        x_reg2[7]) );
  HS65_GS_DFPRQX4 \x_z2_reg[6]  ( .D(n1856), .CP(clk), .RN(rst_n), .Q(x_z2[6])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[6]  ( .D(n1857), .CP(clk), .RN(rst_n), .Q(
        x_reg2[6]) );
  HS65_GS_DFPRQX4 \x_z2_reg[5]  ( .D(n1858), .CP(clk), .RN(rst_n), .Q(x_z2[5])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[5]  ( .D(n1859), .CP(clk), .RN(rst_n), .Q(
        x_reg2[5]) );
  HS65_GS_DFPRQX4 \x_z2_reg[4]  ( .D(n1860), .CP(clk), .RN(rst_n), .Q(x_z2[4])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[4]  ( .D(n1861), .CP(clk), .RN(rst_n), .Q(
        x_reg2[4]) );
  HS65_GS_DFPRQX4 \x_z2_reg[3]  ( .D(n1862), .CP(clk), .RN(rst_n), .Q(x_z2[3])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[3]  ( .D(n1863), .CP(clk), .RN(rst_n), .Q(
        x_reg2[3]) );
  HS65_GS_DFPRQX4 \x_z2_reg[2]  ( .D(n1864), .CP(clk), .RN(rst_n), .Q(x_z2[2])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[2]  ( .D(n1865), .CP(clk), .RN(rst_n), .Q(
        x_reg2[2]) );
  HS65_GS_DFPRQX4 \x_z2_reg[1]  ( .D(n1866), .CP(clk), .RN(rst_n), .Q(x_z2[1])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[1]  ( .D(n1867), .CP(clk), .RN(rst_n), .Q(
        x_reg2[1]) );
  HS65_GS_DFPRQX4 \x_z2_reg[0]  ( .D(n1868), .CP(clk), .RN(rst_n), .Q(x_z2[0])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[0]  ( .D(n1869), .CP(clk), .RN(rst_n), .Q(
        x_reg2[0]) );
  HS65_GS_DFPRQX4 \data_out_reg[15]  ( .D(n1870), .CP(clk), .RN(rst_n), .Q(
        data_out[15]) );
  HS65_GS_DFPRQX4 \y_z1_reg[15]  ( .D(n1871), .CP(clk), .RN(rst_n), .Q(
        y_z1[15]) );
  HS65_GS_DFPRQX4 \y_z2_reg[15]  ( .D(n1872), .CP(clk), .RN(rst_n), .Q(
        y_z2[15]) );
  HS65_GS_DFPRQX4 \data_out_reg[14]  ( .D(n1873), .CP(clk), .RN(rst_n), .Q(
        data_out[14]) );
  HS65_GS_DFPRQX4 \y_z1_reg[14]  ( .D(n1874), .CP(clk), .RN(rst_n), .Q(
        y_z1[14]) );
  HS65_GS_DFPRQX4 \y_z2_reg[14]  ( .D(n1875), .CP(clk), .RN(rst_n), .Q(
        y_z2[14]) );
  HS65_GS_DFPRQX4 \data_out_reg[13]  ( .D(n1876), .CP(clk), .RN(rst_n), .Q(
        data_out[13]) );
  HS65_GS_DFPRQX4 \y_z1_reg[13]  ( .D(n1877), .CP(clk), .RN(rst_n), .Q(
        y_z1[13]) );
  HS65_GS_DFPRQX4 \y_z2_reg[13]  ( .D(n1878), .CP(clk), .RN(rst_n), .Q(
        y_z2[13]) );
  HS65_GS_DFPRQX4 \data_out_reg[12]  ( .D(n1879), .CP(clk), .RN(rst_n), .Q(
        data_out[12]) );
  HS65_GS_DFPRQX4 \y_z1_reg[12]  ( .D(n1880), .CP(clk), .RN(rst_n), .Q(
        y_z1[12]) );
  HS65_GS_DFPRQX4 \y_z2_reg[12]  ( .D(n1881), .CP(clk), .RN(rst_n), .Q(
        y_z2[12]) );
  HS65_GS_DFPRQX4 \data_out_reg[11]  ( .D(n1882), .CP(clk), .RN(rst_n), .Q(
        data_out[11]) );
  HS65_GS_DFPRQX4 \y_z1_reg[11]  ( .D(n1883), .CP(clk), .RN(rst_n), .Q(
        y_z1[11]) );
  HS65_GS_DFPRQX4 \y_z2_reg[11]  ( .D(n1884), .CP(clk), .RN(rst_n), .Q(
        y_z2[11]) );
  HS65_GS_DFPRQX4 \data_out_reg[10]  ( .D(n1885), .CP(clk), .RN(rst_n), .Q(
        data_out[10]) );
  HS65_GS_DFPRQX4 \y_z1_reg[10]  ( .D(n1886), .CP(clk), .RN(rst_n), .Q(
        y_z1[10]) );
  HS65_GS_DFPRQX4 \y_z2_reg[10]  ( .D(n1887), .CP(clk), .RN(rst_n), .Q(
        y_z2[10]) );
  HS65_GS_DFPRQX4 \data_out_reg[9]  ( .D(n1888), .CP(clk), .RN(rst_n), .Q(
        data_out[9]) );
  HS65_GS_DFPRQX4 \y_z1_reg[9]  ( .D(n1889), .CP(clk), .RN(rst_n), .Q(y_z1[9])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[9]  ( .D(n1890), .CP(clk), .RN(rst_n), .Q(y_z2[9])
         );
  HS65_GS_DFPRQX4 \data_out_reg[8]  ( .D(n1891), .CP(clk), .RN(rst_n), .Q(
        data_out[8]) );
  HS65_GS_DFPRQX4 \y_z1_reg[8]  ( .D(n1892), .CP(clk), .RN(rst_n), .Q(y_z1[8])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[8]  ( .D(n1893), .CP(clk), .RN(rst_n), .Q(y_z2[8])
         );
  HS65_GS_DFPRQX4 \data_out_reg[7]  ( .D(n1894), .CP(clk), .RN(rst_n), .Q(
        data_out[7]) );
  HS65_GS_DFPRQX4 \y_z1_reg[7]  ( .D(n1895), .CP(clk), .RN(rst_n), .Q(y_z1[7])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[7]  ( .D(n1896), .CP(clk), .RN(rst_n), .Q(y_z2[7])
         );
  HS65_GS_DFPRQX4 \data_out_reg[6]  ( .D(n1897), .CP(clk), .RN(rst_n), .Q(
        data_out[6]) );
  HS65_GS_DFPRQX4 \y_z1_reg[6]  ( .D(n1898), .CP(clk), .RN(rst_n), .Q(y_z1[6])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[6]  ( .D(n1899), .CP(clk), .RN(rst_n), .Q(y_z2[6])
         );
  HS65_GS_DFPRQX4 \data_out_reg[5]  ( .D(n1900), .CP(clk), .RN(rst_n), .Q(
        data_out[5]) );
  HS65_GS_DFPRQX4 \y_z1_reg[5]  ( .D(n1901), .CP(clk), .RN(rst_n), .Q(y_z1[5])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[5]  ( .D(n1902), .CP(clk), .RN(rst_n), .Q(y_z2[5])
         );
  HS65_GS_DFPRQX4 \data_out_reg[4]  ( .D(n1903), .CP(clk), .RN(rst_n), .Q(
        data_out[4]) );
  HS65_GS_DFPRQX4 \y_z1_reg[4]  ( .D(n1904), .CP(clk), .RN(rst_n), .Q(y_z1[4])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[4]  ( .D(n1905), .CP(clk), .RN(rst_n), .Q(y_z2[4])
         );
  HS65_GS_DFPRQX4 \data_out_reg[3]  ( .D(n1906), .CP(clk), .RN(rst_n), .Q(
        data_out[3]) );
  HS65_GS_DFPRQX4 \y_z1_reg[3]  ( .D(n1907), .CP(clk), .RN(rst_n), .Q(y_z1[3])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[3]  ( .D(n1908), .CP(clk), .RN(rst_n), .Q(y_z2[3])
         );
  HS65_GS_DFPRQX4 \data_out_reg[2]  ( .D(n1909), .CP(clk), .RN(rst_n), .Q(
        data_out[2]) );
  HS65_GS_DFPRQX4 \y_z1_reg[2]  ( .D(n1910), .CP(clk), .RN(rst_n), .Q(y_z1[2])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[2]  ( .D(n1911), .CP(clk), .RN(rst_n), .Q(y_z2[2])
         );
  HS65_GS_DFPRQX4 \data_out_reg[1]  ( .D(n1912), .CP(clk), .RN(rst_n), .Q(
        data_out[1]) );
  HS65_GS_DFPRQX4 \y_z1_reg[1]  ( .D(n1913), .CP(clk), .RN(rst_n), .Q(y_z1[1])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[1]  ( .D(n1914), .CP(clk), .RN(rst_n), .Q(y_z2[1])
         );
  HS65_GS_DFPRQX4 \data_out_reg[0]  ( .D(n1915), .CP(clk), .RN(rst_n), .Q(
        data_out[0]) );
  HS65_GS_DFPRQX4 \y_z1_reg[0]  ( .D(n1916), .CP(clk), .RN(rst_n), .Q(
        \mul_a1/fa1_s1[7] ) );
  HS65_GS_DFPRQX4 \y_z2_reg[0]  ( .D(n1917), .CP(clk), .RN(rst_n), .Q(y_z2[0])
         );
  HS65_GS_NOR2X3 U3 ( .A(\DP_OP_331J1_157_5454/n87 ), .B(n1225), .Z(n1) );
  HS65_GS_AND2X4 U4 ( .A(\mul_b0/fa1_s1_r[29] ), .B(\mul_b0/fa1_s0_r[29] ), 
        .Z(n74) );
  HS65_GSS_XOR2X3 U5 ( .A(\mul_b0/fa1_s0_r[30] ), .B(\mul_b0/fa1_s1_r[30] ), 
        .Z(n73) );
  HS65_GSS_XOR2X3 U6 ( .A(\mul_b0/fa1_s0_r[29] ), .B(\mul_b0/fa1_s1_r[29] ), 
        .Z(n3) );
  HS65_GS_AND2X4 U7 ( .A(\mul_b0/fa1_s0_r[28] ), .B(\mul_b0/fa1_s1_r[28] ), 
        .Z(n2) );
  HS65_GS_FA1X4 U8 ( .A0(\mul_b0/fa1_s2_r[29] ), .B0(n3), .CI(n2), .CO(n617), 
        .S0(n621) );
  HS65_GSS_XOR2X3 U9 ( .A(\mul_b0/fa1_s0_r[28] ), .B(\mul_b0/fa1_s1_r[28] ), 
        .Z(n71) );
  HS65_GS_AND2X4 U10 ( .A(\mul_b0/fa1_s1_r[27] ), .B(\mul_b0/fa1_s0_r[27] ), 
        .Z(n70) );
  HS65_GS_AND2X4 U11 ( .A(\mul_b0/fa1_s0_r[25] ), .B(\mul_b0/fa1_s1_r[25] ), 
        .Z(n5) );
  HS65_GSS_XOR2X3 U12 ( .A(\mul_b0/fa1_s0_r[26] ), .B(\mul_b0/fa1_s1_r[26] ), 
        .Z(n4) );
  HS65_GS_AND2X4 U13 ( .A(\mul_b0/fa1_s1_r[26] ), .B(\mul_b0/fa1_s0_r[26] ), 
        .Z(n69) );
  HS65_GSS_XOR2X3 U14 ( .A(\mul_b0/fa1_s0_r[27] ), .B(\mul_b0/fa1_s1_r[27] ), 
        .Z(n68) );
  HS65_GS_AND2X4 U15 ( .A(\mul_b0/fa1_s0_r[24] ), .B(\mul_b0/fa1_s1_r[24] ), 
        .Z(n63) );
  HS65_GSS_XOR2X3 U16 ( .A(\mul_b0/fa1_s0_r[25] ), .B(\mul_b0/fa1_s1_r[25] ), 
        .Z(n62) );
  HS65_GS_FA1X4 U17 ( .A0(\mul_b0/fa1_s2_r[26] ), .B0(n5), .CI(n4), .CO(n1140), 
        .S0(n1143) );
  HS65_GS_FA1X4 U18 ( .A0(\mul_b0/fa1_s0_r[20] ), .B0(\mul_b0/fa1_s1_r[20] ), 
        .CI(\mul_b0/fa1_c0_r[19] ), .CO(n57), .S0(n6) );
  HS65_GS_FA1X4 U19 ( .A0(\mul_b0/fa1_s0_r[19] ), .B0(\mul_b0/fa1_s1_r[19] ), 
        .CI(\mul_b0/fa1_c0_r[18] ), .CO(n7), .S0(n49) );
  HS65_GS_FA1X4 U20 ( .A0(\mul_b0/fa1_s2_r[20] ), .B0(n7), .CI(n6), .CO(n1160), 
        .S0(n1163) );
  HS65_GS_FA1X4 U21 ( .A0(\mul_b0/fa1_s0_r[17] ), .B0(\mul_b0/fa1_s1_r[17] ), 
        .CI(\mul_b0/fa1_c0_r[16] ), .CO(n52), .S0(n9) );
  HS65_GS_FA1X4 U22 ( .A0(\mul_b0/fa1_s0_r[18] ), .B0(\mul_b0/fa1_s1_r[18] ), 
        .CI(\mul_b0/fa1_c0_r[17] ), .CO(n50), .S0(n51) );
  HS65_GS_FA1X4 U23 ( .A0(\mul_b0/fa1_s2_r[17] ), .B0(n9), .CI(n8), .CO(n638), 
        .S0(n47) );
  HS65_GS_FA1X4 U24 ( .A0(\mul_b0/fa1_s0_r[16] ), .B0(\mul_b0/fa1_s1_r[16] ), 
        .CI(\mul_b0/fa1_c0_r[15] ), .CO(n8), .S0(n41) );
  HS65_GS_NAND2X2 U25 ( .A(n47), .B(n46), .Z(n48) );
  HS65_GS_FA1X4 U26 ( .A0(\mul_b0/fa1_s0_r[15] ), .B0(\mul_b0/fa1_s1_r[15] ), 
        .CI(\mul_b0/fa1_c0_r[14] ), .CO(n42), .S0(n43) );
  HS65_GS_FA1X4 U27 ( .A0(\mul_b0/fa1_s0_r[14] ), .B0(\mul_b0/fa1_s1_r[14] ), 
        .CI(\mul_b0/fa1_c0_r[13] ), .CO(n44), .S0(n10) );
  HS65_GS_FA1X4 U28 ( .A0(\mul_b0/fa1_s2_r[14] ), .B0(n11), .CI(n10), .CO(n39), 
        .S0(n37) );
  HS65_GS_FA1X4 U29 ( .A0(\mul_b0/fa1_s0_r[13] ), .B0(\mul_b0/fa1_s1_r[13] ), 
        .CI(\mul_b0/fa1_c0_r[12] ), .CO(n11), .S0(n13) );
  HS65_GS_NAND2X2 U30 ( .A(n37), .B(n36), .Z(n38) );
  HS65_GS_NAND2X2 U31 ( .A(n40), .B(n39), .Z(n12) );
  HS65_GS_OAI21X2 U32 ( .A(n40), .B(n39), .C(n12), .Z(n1801) );
  HS65_GS_NAND2X2 U33 ( .A(n38), .B(n1801), .Z(n1803) );
  HS65_GS_FA1X4 U34 ( .A0(\mul_b0/fa1_s2_r[13] ), .B0(n14), .CI(n13), .CO(n36), 
        .S0(n35) );
  HS65_GS_FA1X4 U35 ( .A0(\mul_b0/fa1_s0_r[12] ), .B0(\mul_b0/fa1_s1_r[12] ), 
        .CI(\mul_b0/fa1_c0_r[11] ), .CO(n14), .S0(n15) );
  HS65_GS_FA1X4 U36 ( .A0(\mul_b0/fa1_s2_r[12] ), .B0(n16), .CI(n15), .CO(n34), 
        .S0(n32) );
  HS65_GS_FA1X4 U37 ( .A0(\mul_b0/fa1_s0_r[11] ), .B0(\mul_b0/fa1_s1_r[11] ), 
        .CI(\mul_b0/fa1_c0_r[10] ), .CO(n16), .S0(n29) );
  HS65_GS_FA1X4 U38 ( .A0(\mul_b0/fa1_s0_r[10] ), .B0(\mul_b0/fa1_s1_r[10] ), 
        .CI(\mul_b0/fa1_c0_r[9] ), .CO(n30), .S0(n26) );
  HS65_GS_NOR2X2 U39 ( .A(n27), .B(n26), .Z(n24) );
  HS65_GS_FA1X4 U40 ( .A0(\mul_b0/fa1_s0_r[8] ), .B0(\mul_b0/fa1_s1_r[8] ), 
        .CI(\mul_b0/fa1_c0_r[7] ), .CO(n22), .S0(n19) );
  HS65_GS_AND2X4 U41 ( .A(\mul_b0/fa1_c0_r[5] ), .B(\mul_b0/fa1_s0_r[6] ), .Z(
        n17) );
  HS65_GS_PAOI2X1 U42 ( .A(\mul_b0/fa1_s0_r[7] ), .B(\mul_b0/fa1_c0_r[6] ), 
        .P(n17), .Z(n18) );
  HS65_GS_NOR2AX3 U43 ( .A(n19), .B(n18), .Z(n21) );
  HS65_GS_FA1X4 U44 ( .A0(\mul_b0/fa1_s0_r[9] ), .B0(\mul_b0/fa1_s1_r[9] ), 
        .CI(\mul_b0/fa1_c0_r[8] ), .CO(n27), .S0(n20) );
  HS65_GS_PAOI2X1 U45 ( .A(n22), .B(n21), .P(n20), .Z(n23) );
  HS65_GS_NOR2X2 U46 ( .A(n24), .B(n23), .Z(n25) );
  HS65_GS_AO12X4 U47 ( .A(n27), .B(n26), .C(n25), .Z(n28) );
  HS65_GS_PAOI2X1 U48 ( .A(n30), .B(n29), .P(n28), .Z(n31) );
  HS65_GS_NOR2AX3 U49 ( .A(n32), .B(n31), .Z(n33) );
  HS65_GS_PAO2X4 U50 ( .A(n35), .B(n34), .P(n33), .Z(n1173) );
  HS65_GSS_XOR2X3 U51 ( .A(n37), .B(n36), .Z(n1172) );
  HS65_GS_NAND2X2 U52 ( .A(n1173), .B(n1172), .Z(n1800) );
  HS65_GS_OAI21X2 U53 ( .A(n1801), .B(n38), .C(n1800), .Z(n1799) );
  HS65_GS_AOI22X1 U54 ( .A(n40), .B(n39), .C(n1803), .D(n1799), .Z(n648) );
  HS65_GS_FA1X4 U55 ( .A0(\mul_b0/fa1_s2_r[16] ), .B0(n42), .CI(n41), .CO(n46), 
        .S0(n646) );
  HS65_GS_FA1X4 U56 ( .A0(\mul_b0/fa1_s2_r[15] ), .B0(n44), .CI(n43), .CO(n645), .S0(n40) );
  HS65_GS_NAND2X2 U57 ( .A(n646), .B(n645), .Z(n644) );
  HS65_GS_NOR2X2 U58 ( .A(n646), .B(n645), .Z(n45) );
  HS65_GS_AOI12X2 U59 ( .A(n648), .B(n644), .C(n45), .Z(n1170) );
  HS65_GSS_XOR2X3 U60 ( .A(n47), .B(n46), .Z(n1169) );
  HS65_GS_NAND2X2 U61 ( .A(n1170), .B(n1169), .Z(n1168) );
  HS65_GS_NAND2X2 U62 ( .A(n48), .B(n1168), .Z(n640) );
  HS65_GS_PAOI2X1 U63 ( .A(n638), .B(n639), .P(n640), .Z(n636) );
  HS65_GS_FA1X4 U64 ( .A0(\mul_b0/fa1_s2_r[19] ), .B0(n50), .CI(n49), .CO(
        n1164), .S0(n54) );
  HS65_GS_FA1X4 U65 ( .A0(\mul_b0/fa1_s2_r[18] ), .B0(n52), .CI(n51), .CO(n53), 
        .S0(n639) );
  HS65_GS_NAND2X2 U66 ( .A(n54), .B(n53), .Z(n55) );
  HS65_GS_OAI21X2 U67 ( .A(n54), .B(n53), .C(n55), .Z(n635) );
  HS65_GS_OAI21X2 U68 ( .A(n636), .B(n635), .C(n55), .Z(n1162) );
  HS65_GS_FA1X4 U69 ( .A0(\mul_b0/fa1_s2_r[21] ), .B0(n57), .CI(n56), .CO(
        n1155), .S0(n1159) );
  HS65_GS_FA1X4 U70 ( .A0(\mul_b0/fa1_s0_r[21] ), .B0(\mul_b0/fa1_s1_r[21] ), 
        .CI(\mul_b0/fa1_c0_r[20] ), .CO(n59), .S0(n56) );
  HS65_GSS_XOR2X3 U71 ( .A(\mul_b0/fa1_s0_r[22] ), .B(\mul_b0/fa1_s1_r[22] ), 
        .Z(n58) );
  HS65_GS_FA1X4 U72 ( .A0(\mul_b0/fa1_s2_r[22] ), .B0(n59), .CI(n58), .CO(
        n1151), .S0(n1154) );
  HS65_GSS_XOR2X3 U73 ( .A(\mul_b0/fa1_s0_r[23] ), .B(\mul_b0/fa1_s1_r[23] ), 
        .Z(n61) );
  HS65_GS_AND2X4 U74 ( .A(\mul_b0/fa1_s1_r[22] ), .B(\mul_b0/fa1_s0_r[22] ), 
        .Z(n60) );
  HS65_GS_FA1X4 U75 ( .A0(\mul_b0/fa1_s2_r[23] ), .B0(n61), .CI(n60), .CO(
        n1147), .S0(n1150) );
  HS65_GS_AND2X4 U76 ( .A(\mul_b0/fa1_s1_r[23] ), .B(\mul_b0/fa1_s0_r[23] ), 
        .Z(n65) );
  HS65_GSS_XOR2X3 U77 ( .A(\mul_b0/fa1_s0_r[24] ), .B(\mul_b0/fa1_s1_r[24] ), 
        .Z(n64) );
  HS65_GS_FA1X4 U78 ( .A0(\mul_b0/fa1_s2_r[25] ), .B0(n63), .CI(n62), .CO(
        n1144), .S0(n67) );
  HS65_GS_FA1X4 U79 ( .A0(\mul_b0/fa1_s2_r[24] ), .B0(n65), .CI(n64), .CO(n66), 
        .S0(n1146) );
  HS65_GSS_XOR2X3 U80 ( .A(n67), .B(n66), .Z(n633) );
  HS65_GS_AO22X4 U81 ( .A(n632), .B(n633), .C(n67), .D(n66), .Z(n1142) );
  HS65_GS_FA1X4 U82 ( .A0(\mul_b0/fa1_s2_r[27] ), .B0(n69), .CI(n68), .CO(
        n1135), .S0(n1139) );
  HS65_GS_FA1X4 U83 ( .A0(\mul_b0/fa1_s2_r[28] ), .B0(n71), .CI(n70), .CO(n620), .S0(n1134) );
  HS65_GS_IVX2 U84 ( .A(n72), .Z(n624) );
  HS65_GSS_XOR2X3 U85 ( .A(\mul_b0/fa1_s0_r[31] ), .B(\mul_b0/fa1_s1_r[31] ), 
        .Z(n79) );
  HS65_GS_AND2X4 U86 ( .A(\mul_b0/fa1_s1_r[30] ), .B(\mul_b0/fa1_s0_r[30] ), 
        .Z(n78) );
  HS65_GS_FA1X4 U87 ( .A0(\mul_b0/fa1_s2_r[30] ), .B0(n74), .CI(n73), .CO(n75), 
        .S0(n618) );
  HS65_GS_NAND2X2 U88 ( .A(n76), .B(n75), .Z(n77) );
  HS65_GS_OAI21X2 U89 ( .A(n76), .B(n75), .C(n77), .Z(n623) );
  HS65_GS_NOR2X2 U90 ( .A(n624), .B(n623), .Z(n622) );
  HS65_GS_IVX2 U91 ( .A(n77), .Z(n82) );
  HS65_GS_AND2X4 U92 ( .A(\mul_b0/fa1_s1_r[31] ), .B(\mul_b0/fa1_s0_r[31] ), 
        .Z(n85) );
  HS65_GSS_XOR2X3 U93 ( .A(\mul_b0/fa1_s0_r[32] ), .B(\mul_b0/fa1_s1_r[32] ), 
        .Z(n84) );
  HS65_GS_FA1X4 U94 ( .A0(\mul_b0/fa1_s2_r[31] ), .B0(n79), .CI(n78), .CO(n80), 
        .S0(n76) );
  HS65_GS_FA1X4 U95 ( .A0(n82), .B0(n81), .CI(n80), .CO(n83), .S0(n615) );
  HS65_GS_AOI12X2 U96 ( .A(n622), .B(n615), .C(n83), .Z(n90) );
  HS65_GS_AND2X4 U97 ( .A(\mul_b0/fa1_s1_r[32] ), .B(\mul_b0/fa1_s0_r[32] ), 
        .Z(n87) );
  HS65_GS_FA1X4 U98 ( .A0(\mul_b0/fa1_s2_r[32] ), .B0(n85), .CI(n84), .CO(n86), 
        .S0(n81) );
  HS65_GSS_XOR3X2 U99 ( .A(n87), .B(n86), .C(\mul_b0/fa1_s2_r[33] ), .Z(n88)
         );
  HS65_GSS_XOR3X2 U100 ( .A(\mul_b0/fa1_s0_r[33] ), .B(\mul_b0/fa1_s1_r[33] ), 
        .C(n88), .Z(n89) );
  HS65_GSS_XNOR2X3 U101 ( .A(n90), .B(n89), .Z(\mul_b0/result_sat[15] ) );
  HS65_GS_AND2X4 U102 ( .A(\mul_a2/fa1_s1_r[28] ), .B(\mul_a2/fa1_s0_r[28] ), 
        .Z(n92) );
  HS65_GSS_XOR2X3 U103 ( .A(\mul_a2/fa1_s0_r[29] ), .B(\mul_a2/fa1_s1_r[29] ), 
        .Z(n91) );
  HS65_GSS_XOR2X3 U104 ( .A(\mul_a2/fa1_s0_r[30] ), .B(\mul_a2/fa1_s1_r[30] ), 
        .Z(n172) );
  HS65_GS_AND2X4 U105 ( .A(\mul_a2/fa1_s1_r[29] ), .B(\mul_a2/fa1_s0_r[29] ), 
        .Z(n171) );
  HS65_GS_AND2X4 U106 ( .A(\mul_a2/fa1_s1_r[27] ), .B(\mul_a2/fa1_s0_r[27] ), 
        .Z(n164) );
  HS65_GSS_XOR2X3 U107 ( .A(\mul_a2/fa1_s0_r[28] ), .B(\mul_a2/fa1_s1_r[28] ), 
        .Z(n163) );
  HS65_GS_FA1X4 U108 ( .A0(\mul_a2/fa1_s2_r[29] ), .B0(n92), .CI(n91), .CO(
        n653), .S0(n655) );
  HS65_GS_AND2X4 U109 ( .A(\mul_a2/fa1_s1_r[21] ), .B(\mul_a2/fa1_s0_r[21] ), 
        .Z(n94) );
  HS65_GSS_XOR2X3 U110 ( .A(\mul_a2/fa1_s1_r[22] ), .B(\mul_a2/fa1_s0_r[22] ), 
        .Z(n93) );
  HS65_GS_AND2X4 U111 ( .A(\mul_a2/fa1_s0_r[22] ), .B(\mul_a2/fa1_s1_r[22] ), 
        .Z(n156) );
  HS65_GSS_XOR2X3 U112 ( .A(\mul_a2/fa1_s1_r[23] ), .B(\mul_a2/fa1_s0_r[23] ), 
        .Z(n155) );
  HS65_GS_AND2X4 U113 ( .A(\mul_a2/fa1_s1_r[20] ), .B(\mul_a2/fa1_s0_r[20] ), 
        .Z(n96) );
  HS65_GSS_XOR2X3 U114 ( .A(\mul_a2/fa1_s0_r[21] ), .B(\mul_a2/fa1_s1_r[21] ), 
        .Z(n95) );
  HS65_GS_FA1X4 U115 ( .A0(\mul_a2/fa1_s2_r[22] ), .B0(n94), .CI(n93), .CO(
        n1326), .S0(n1329) );
  HS65_GSS_XOR2X3 U116 ( .A(\mul_a2/fa1_s0_r[20] ), .B(\mul_a2/fa1_s1_r[20] ), 
        .Z(n98) );
  HS65_GS_AND2X4 U117 ( .A(\mul_a2/fa1_s1_r[19] ), .B(\mul_a2/fa1_s0_r[19] ), 
        .Z(n97) );
  HS65_GS_FA1X4 U118 ( .A0(\mul_a2/fa1_s2_r[21] ), .B0(n96), .CI(n95), .CO(
        n1330), .S0(n1333) );
  HS65_GS_AND2X4 U119 ( .A(\mul_a2/fa1_s1_r[18] ), .B(\mul_a2/fa1_s0_r[18] ), 
        .Z(n149) );
  HS65_GSS_XOR2X3 U120 ( .A(\mul_a2/fa1_s0_r[19] ), .B(\mul_a2/fa1_s1_r[19] ), 
        .Z(n148) );
  HS65_GS_FA1X4 U121 ( .A0(\mul_a2/fa1_s2_r[20] ), .B0(n98), .CI(n97), .CO(
        n1334), .S0(n1337) );
  HS65_GS_PAO2X4 U122 ( .A(\mul_a2/fa1_c0_r[16] ), .B(\mul_a2/fa1_s1_r[17] ), 
        .P(\mul_a2/fa1_s0_r[17] ), .Z(n151) );
  HS65_GSS_XOR2X3 U123 ( .A(\mul_a2/fa1_s0_r[18] ), .B(\mul_a2/fa1_s1_r[18] ), 
        .Z(n150) );
  HS65_GS_PAO2X4 U124 ( .A(\mul_a2/fa1_s1_r[16] ), .B(\mul_a2/fa1_s0_r[16] ), 
        .P(\mul_a2/fa1_c0_r[15] ), .Z(n100) );
  HS65_GSS_XOR3X2 U125 ( .A(\mul_a2/fa1_c0_r[16] ), .B(\mul_a2/fa1_s1_r[17] ), 
        .C(\mul_a2/fa1_s0_r[17] ), .Z(n99) );
  HS65_GS_FA1X4 U126 ( .A0(\mul_a2/fa1_s2_r[17] ), .B0(n100), .CI(n99), .CO(
        n679), .S0(n146) );
  HS65_GS_PAO2X4 U127 ( .A(\mul_a2/fa1_c0_r[14] ), .B(\mul_a2/fa1_s1_r[15] ), 
        .P(\mul_a2/fa1_s0_r[15] ), .Z(n143) );
  HS65_GSS_XOR3X2 U128 ( .A(\mul_a2/fa1_s1_r[16] ), .B(\mul_a2/fa1_s0_r[16] ), 
        .C(\mul_a2/fa1_c0_r[15] ), .Z(n142) );
  HS65_GS_NAND2X2 U129 ( .A(n146), .B(n145), .Z(n147) );
  HS65_GS_PAO2X4 U130 ( .A(\mul_a2/fa1_c0_r[13] ), .B(\mul_a2/fa1_s1_r[14] ), 
        .P(\mul_a2/fa1_s0_r[14] ), .Z(n141) );
  HS65_GSS_XOR3X2 U131 ( .A(\mul_a2/fa1_c0_r[14] ), .B(\mul_a2/fa1_s1_r[15] ), 
        .C(\mul_a2/fa1_s0_r[15] ), .Z(n140) );
  HS65_GS_PAO2X4 U132 ( .A(\mul_a2/fa1_c0_r[12] ), .B(\mul_a2/fa1_s1_r[13] ), 
        .P(\mul_a2/fa1_s0_r[13] ), .Z(n102) );
  HS65_GSS_XOR3X2 U133 ( .A(\mul_a2/fa1_c0_r[13] ), .B(\mul_a2/fa1_s1_r[14] ), 
        .C(\mul_a2/fa1_s0_r[14] ), .Z(n101) );
  HS65_GSS_XOR3X2 U134 ( .A(\mul_a2/fa1_c0_r[12] ), .B(\mul_a2/fa1_s1_r[13] ), 
        .C(\mul_a2/fa1_s0_r[13] ), .Z(n105) );
  HS65_GS_PAO2X4 U135 ( .A(\mul_a2/fa1_s1_r[12] ), .B(\mul_a2/fa1_s0_r[12] ), 
        .P(\mul_a2/fa1_c0_r[11] ), .Z(n104) );
  HS65_GS_PAOI2X1 U136 ( .A(n105), .B(n104), .P(\mul_a2/fa1_s2_r[13] ), .Z(
        n136) );
  HS65_GS_FA1X4 U137 ( .A0(\mul_a2/fa1_s2_r[14] ), .B0(n102), .CI(n101), .CO(
        n138), .S0(n135) );
  HS65_GS_NAND2AX4 U138 ( .A(n136), .B(n135), .Z(n137) );
  HS65_GS_NAND2X2 U139 ( .A(n139), .B(n138), .Z(n103) );
  HS65_GS_OAI21X2 U140 ( .A(n139), .B(n138), .C(n103), .Z(n1758) );
  HS65_GS_NAND2X2 U141 ( .A(n137), .B(n1758), .Z(n1760) );
  HS65_GSS_XOR2X3 U142 ( .A(n105), .B(n104), .Z(n134) );
  HS65_GS_PAO2X4 U143 ( .A(\mul_a2/fa1_c0_r[10] ), .B(\mul_a2/fa1_s1_r[11] ), 
        .P(\mul_a2/fa1_s0_r[11] ), .Z(n131) );
  HS65_GSS_XOR3X2 U144 ( .A(\mul_a2/fa1_s1_r[12] ), .B(\mul_a2/fa1_s0_r[12] ), 
        .C(\mul_a2/fa1_c0_r[11] ), .Z(n130) );
  HS65_GS_AND2X4 U145 ( .A(\mul_a2/fa1_c0_r[8] ), .B(\mul_a2/fa1_s0_r[9] ), 
        .Z(n125) );
  HS65_GSS_XOR2X3 U146 ( .A(\mul_a2/fa1_c0_r[9] ), .B(\mul_a2/fa1_s0_r[10] ), 
        .Z(n124) );
  HS65_GS_AND2X4 U147 ( .A(\mul_a2/fa1_c0_r[6] ), .B(\mul_a2/fa1_s0_r[7] ), 
        .Z(n119) );
  HS65_GSS_XOR2X3 U148 ( .A(\mul_a2/fa1_c0_r[7] ), .B(\mul_a2/fa1_s0_r[8] ), 
        .Z(n118) );
  HS65_GS_AND2X4 U149 ( .A(\mul_a2/fa1_c0_r[4] ), .B(\mul_a2/fa1_s0_r[5] ), 
        .Z(n113) );
  HS65_GSS_XOR2X3 U150 ( .A(\mul_a2/fa1_c0_r[5] ), .B(\mul_a2/fa1_s0_r[6] ), 
        .Z(n112) );
  HS65_GSS_XOR2X3 U151 ( .A(\mul_a2/fa1_c0_r[4] ), .B(\mul_a2/fa1_s0_r[5] ), 
        .Z(n110) );
  HS65_GS_AND2X4 U152 ( .A(\mul_a2/fa1_c0_r[3] ), .B(\mul_a2/fa1_s0_r[4] ), 
        .Z(n109) );
  HS65_GS_NAND2X2 U153 ( .A(\mul_a2/fa1_c0_r[2] ), .B(\mul_a2/fa1_s0_r[3] ), 
        .Z(n107) );
  HS65_GSS_XNOR2X3 U154 ( .A(\mul_a2/fa1_c0_r[3] ), .B(\mul_a2/fa1_s0_r[4] ), 
        .Z(n106) );
  HS65_GS_NOR2X2 U155 ( .A(n107), .B(n106), .Z(n108) );
  HS65_GS_PAO2X4 U156 ( .A(n110), .B(n109), .P(n108), .Z(n111) );
  HS65_GS_PAO2X4 U157 ( .A(n113), .B(n112), .P(n111), .Z(n116) );
  HS65_GS_AND2X4 U158 ( .A(\mul_a2/fa1_c0_r[5] ), .B(\mul_a2/fa1_s0_r[6] ), 
        .Z(n115) );
  HS65_GSS_XOR2X3 U159 ( .A(\mul_a2/fa1_c0_r[6] ), .B(\mul_a2/fa1_s0_r[7] ), 
        .Z(n114) );
  HS65_GS_PAO2X4 U160 ( .A(n116), .B(n115), .P(n114), .Z(n117) );
  HS65_GS_PAO2X4 U161 ( .A(n119), .B(n118), .P(n117), .Z(n122) );
  HS65_GS_AND2X4 U162 ( .A(\mul_a2/fa1_c0_r[7] ), .B(\mul_a2/fa1_s0_r[8] ), 
        .Z(n121) );
  HS65_GSS_XOR2X3 U163 ( .A(\mul_a2/fa1_c0_r[8] ), .B(\mul_a2/fa1_s0_r[9] ), 
        .Z(n120) );
  HS65_GS_PAO2X4 U164 ( .A(n122), .B(n121), .P(n120), .Z(n123) );
  HS65_GS_PAO2X4 U165 ( .A(n125), .B(n124), .P(n123), .Z(n128) );
  HS65_GSS_XOR3X2 U166 ( .A(\mul_a2/fa1_c0_r[10] ), .B(\mul_a2/fa1_s1_r[11] ), 
        .C(\mul_a2/fa1_s0_r[11] ), .Z(n127) );
  HS65_GS_AND2X4 U167 ( .A(\mul_a2/fa1_c0_r[9] ), .B(\mul_a2/fa1_s0_r[10] ), 
        .Z(n126) );
  HS65_GS_PAO2X4 U168 ( .A(n128), .B(n127), .P(n126), .Z(n129) );
  HS65_GS_PAOI2X1 U169 ( .A(n131), .B(n130), .P(n129), .Z(n133) );
  HS65_GS_NOR2X2 U170 ( .A(n134), .B(\mul_a2/fa1_s2_r[13] ), .Z(n132) );
  HS65_GS_AOI112X2 U171 ( .A(n134), .B(\mul_a2/fa1_s2_r[13] ), .C(n133), .D(
        n132), .Z(n1347) );
  HS65_GSS_XNOR2X3 U172 ( .A(n136), .B(n135), .Z(n1346) );
  HS65_GS_NAND2X2 U173 ( .A(n1347), .B(n1346), .Z(n1757) );
  HS65_GS_OAI21X2 U174 ( .A(n1758), .B(n137), .C(n1757), .Z(n1756) );
  HS65_GS_AOI22X1 U175 ( .A(n139), .B(n138), .C(n1760), .D(n1756), .Z(n688) );
  HS65_GS_FA1X4 U176 ( .A0(\mul_a2/fa1_s2_r[15] ), .B0(n141), .CI(n140), .CO(
        n686), .S0(n139) );
  HS65_GS_FA1X4 U177 ( .A0(\mul_a2/fa1_s2_r[16] ), .B0(n143), .CI(n142), .CO(
        n145), .S0(n685) );
  HS65_GS_NAND2X2 U178 ( .A(n686), .B(n685), .Z(n684) );
  HS65_GS_NOR2X2 U179 ( .A(n686), .B(n685), .Z(n144) );
  HS65_GS_AOI12X2 U180 ( .A(n688), .B(n684), .C(n144), .Z(n1344) );
  HS65_GSS_XOR2X3 U181 ( .A(n146), .B(n145), .Z(n1343) );
  HS65_GS_NAND2X2 U182 ( .A(n1344), .B(n1343), .Z(n1342) );
  HS65_GS_NAND2X2 U183 ( .A(n147), .B(n1342), .Z(n680) );
  HS65_GS_PAOI2X1 U184 ( .A(n678), .B(n679), .P(n680), .Z(n676) );
  HS65_GS_FA1X4 U185 ( .A0(\mul_a2/fa1_s2_r[19] ), .B0(n149), .CI(n148), .CO(
        n1338), .S0(n153) );
  HS65_GS_FA1X4 U186 ( .A0(\mul_a2/fa1_s2_r[18] ), .B0(n151), .CI(n150), .CO(
        n152), .S0(n678) );
  HS65_GS_NAND2X2 U187 ( .A(n153), .B(n152), .Z(n154) );
  HS65_GS_OAI21X2 U188 ( .A(n153), .B(n152), .C(n154), .Z(n675) );
  HS65_GS_OAI21X2 U189 ( .A(n676), .B(n675), .C(n154), .Z(n1336) );
  HS65_GS_FA1X4 U190 ( .A0(\mul_a2/fa1_s2_r[23] ), .B0(n156), .CI(n155), .CO(
        n1321), .S0(n1325) );
  HS65_GS_AND2X4 U191 ( .A(\mul_a2/fa1_s0_r[23] ), .B(\mul_a2/fa1_s1_r[23] ), 
        .Z(n158) );
  HS65_GSS_XOR2X3 U192 ( .A(\mul_a2/fa1_s1_r[24] ), .B(\mul_a2/fa1_s0_r[24] ), 
        .Z(n157) );
  HS65_GS_FA1X4 U193 ( .A0(\mul_a2/fa1_s2_r[24] ), .B0(n158), .CI(n157), .CO(
        n1317), .S0(n1320) );
  HS65_GSS_XOR2X3 U194 ( .A(\mul_a2/fa1_s1_r[25] ), .B(\mul_a2/fa1_s0_r[25] ), 
        .Z(n160) );
  HS65_GS_AND2X4 U195 ( .A(\mul_a2/fa1_s0_r[24] ), .B(\mul_a2/fa1_s1_r[24] ), 
        .Z(n159) );
  HS65_GS_FA1X4 U196 ( .A0(\mul_a2/fa1_s2_r[25] ), .B0(n160), .CI(n159), .CO(
        n1313), .S0(n1316) );
  HS65_GSS_XOR2X3 U197 ( .A(\mul_a2/fa1_s1_r[26] ), .B(\mul_a2/fa1_s0_r[26] ), 
        .Z(n162) );
  HS65_GS_AND2X4 U198 ( .A(\mul_a2/fa1_s0_r[25] ), .B(\mul_a2/fa1_s1_r[25] ), 
        .Z(n161) );
  HS65_GS_AND2X4 U199 ( .A(\mul_a2/fa1_s0_r[26] ), .B(\mul_a2/fa1_s1_r[26] ), 
        .Z(n166) );
  HS65_GSS_XOR2X3 U200 ( .A(\mul_a2/fa1_s0_r[27] ), .B(\mul_a2/fa1_s1_r[27] ), 
        .Z(n165) );
  HS65_GS_FA1X4 U201 ( .A0(\mul_a2/fa1_s2_r[26] ), .B0(n162), .CI(n161), .CO(
        n669), .S0(n1312) );
  HS65_GS_PAOI2X1 U202 ( .A(n672), .B(n670), .P(n669), .Z(n667) );
  HS65_GS_FA1X4 U203 ( .A0(\mul_a2/fa1_s2_r[28] ), .B0(n164), .CI(n163), .CO(
        n656), .S0(n168) );
  HS65_GS_FA1X4 U204 ( .A0(\mul_a2/fa1_s2_r[27] ), .B0(n166), .CI(n165), .CO(
        n167), .S0(n670) );
  HS65_GS_NAND2X2 U205 ( .A(n168), .B(n167), .Z(n169) );
  HS65_GS_OAI21X2 U206 ( .A(n168), .B(n167), .C(n169), .Z(n668) );
  HS65_GS_OAI21X2 U207 ( .A(n667), .B(n668), .C(n169), .Z(n654) );
  HS65_GS_IVX2 U208 ( .A(n170), .Z(n659) );
  HS65_GSS_XOR2X3 U209 ( .A(\mul_a2/fa1_s1_r[31] ), .B(\mul_a2/fa1_s0_r[31] ), 
        .Z(n177) );
  HS65_GS_AND2X4 U210 ( .A(\mul_a2/fa1_s1_r[30] ), .B(\mul_a2/fa1_s0_r[30] ), 
        .Z(n176) );
  HS65_GS_FA1X4 U211 ( .A0(\mul_a2/fa1_s2_r[30] ), .B0(n172), .CI(n171), .CO(
        n173), .S0(n652) );
  HS65_GS_NAND2X2 U212 ( .A(n174), .B(n173), .Z(n175) );
  HS65_GS_OAI21X2 U213 ( .A(n174), .B(n173), .C(n175), .Z(n658) );
  HS65_GS_NOR2X2 U214 ( .A(n659), .B(n658), .Z(n657) );
  HS65_GS_IVX2 U215 ( .A(n175), .Z(n180) );
  HS65_GS_FA1X4 U216 ( .A0(\mul_a2/fa1_s2_r[31] ), .B0(n177), .CI(n176), .CO(
        n179), .S0(n174) );
  HS65_GSS_XOR2X3 U217 ( .A(\mul_a2/fa1_s1_r[32] ), .B(\mul_a2/fa1_s0_r[32] ), 
        .Z(n183) );
  HS65_GS_AND2X4 U218 ( .A(\mul_a2/fa1_s0_r[31] ), .B(\mul_a2/fa1_s1_r[31] ), 
        .Z(n182) );
  HS65_GS_FA1X4 U219 ( .A0(n180), .B0(n179), .CI(n178), .CO(n181), .S0(n650)
         );
  HS65_GS_AOI12X2 U220 ( .A(n657), .B(n650), .C(n181), .Z(n188) );
  HS65_GS_FA1X4 U221 ( .A0(\mul_a2/fa1_s2_r[32] ), .B0(n183), .CI(n182), .CO(
        n186), .S0(n178) );
  HS65_GS_NAND2X2 U222 ( .A(\mul_a2/fa1_s1_r[32] ), .B(\mul_a2/fa1_s0_r[32] ), 
        .Z(n184) );
  HS65_GSS_XNOR3X2 U223 ( .A(n184), .B(\mul_a2/fa1_s0_r[33] ), .C(
        \mul_a2/fa1_s1_r[33] ), .Z(n185) );
  HS65_GSS_XOR3X2 U224 ( .A(\mul_a2/fa1_s2_r[33] ), .B(n186), .C(n185), .Z(
        n187) );
  HS65_GSS_XNOR2X3 U225 ( .A(n188), .B(n187), .Z(\mul_a2/result_sat[15] ) );
  HS65_GS_BFX4 U226 ( .A(valid_in), .Z(n1821) );
  HS65_GS_IVX2 U227 ( .A(x_z1[15]), .Z(n1438) );
  HS65_GS_PAO2X4 U228 ( .A(\mul_b2/fa1_c0_r[31] ), .B(\mul_b2/fa1_s1_r[32] ), 
        .P(\mul_b2/fa1_s0_r[32] ), .Z(n409) );
  HS65_GSS_XOR3X2 U229 ( .A(\mul_b2/fa1_c0_r[31] ), .B(\mul_b2/fa1_s1_r[32] ), 
        .C(\mul_b2/fa1_s0_r[32] ), .Z(n190) );
  HS65_GS_PAO2X4 U230 ( .A(\mul_b2/fa1_c0_r[30] ), .B(\mul_b2/fa1_s1_r[31] ), 
        .P(\mul_b2/fa1_s0_r[31] ), .Z(n189) );
  HS65_GS_FA1X4 U231 ( .A0(n190), .B0(\mul_b2/fa1_s2_r[32] ), .CI(n189), .CO(
        n405), .S0(n191) );
  HS65_GSS_XOR3X2 U232 ( .A(\mul_b2/fa1_c0_r[30] ), .B(\mul_b2/fa1_s1_r[31] ), 
        .C(\mul_b2/fa1_s0_r[31] ), .Z(n399) );
  HS65_GS_PAO2X4 U233 ( .A(\mul_b2/fa1_c0_r[29] ), .B(\mul_b2/fa1_s1_r[30] ), 
        .P(\mul_b2/fa1_s0_r[30] ), .Z(n398) );
  HS65_GS_AND2X4 U234 ( .A(n191), .B(n192), .Z(n403) );
  HS65_GSS_XNOR2X3 U235 ( .A(n192), .B(n191), .Z(n830) );
  HS65_GSS_XOR3X2 U236 ( .A(\mul_b2/fa1_c0_r[28] ), .B(\mul_b2/fa1_s1_r[29] ), 
        .C(\mul_b2/fa1_s0_r[29] ), .Z(n195) );
  HS65_GS_PAO2X4 U237 ( .A(\mul_b2/fa1_c0_r[27] ), .B(\mul_b2/fa1_s1_r[28] ), 
        .P(\mul_b2/fa1_s0_r[28] ), .Z(n194) );
  HS65_GS_PAO2X4 U238 ( .A(\mul_b2/fa1_c0_r[28] ), .B(\mul_b2/fa1_s1_r[29] ), 
        .P(\mul_b2/fa1_s0_r[29] ), .Z(n397) );
  HS65_GSS_XOR3X2 U239 ( .A(\mul_b2/fa1_c0_r[29] ), .B(\mul_b2/fa1_s1_r[30] ), 
        .C(\mul_b2/fa1_s0_r[30] ), .Z(n396) );
  HS65_GS_IVX2 U240 ( .A(n395), .Z(n394) );
  HS65_GS_NAND2X2 U241 ( .A(n393), .B(n395), .Z(n824) );
  HS65_GS_PAO2X4 U242 ( .A(\mul_b2/fa1_s1_r[27] ), .B(\mul_b2/fa1_s0_r[27] ), 
        .P(\mul_b2/fa1_c0_r[26] ), .Z(n193) );
  HS65_GSS_XOR2X3 U243 ( .A(n193), .B(\mul_b2/fa1_s2_r[28] ), .Z(n388) );
  HS65_GSS_XOR3X2 U244 ( .A(\mul_b2/fa1_c0_r[27] ), .B(\mul_b2/fa1_s1_r[28] ), 
        .C(\mul_b2/fa1_s0_r[28] ), .Z(n389) );
  HS65_GS_NAND2X2 U245 ( .A(n388), .B(n389), .Z(n380) );
  HS65_GS_IVX2 U246 ( .A(n380), .Z(n196) );
  HS65_GS_AND2X4 U247 ( .A(n193), .B(\mul_b2/fa1_s2_r[28] ), .Z(n387) );
  HS65_GS_FA1X4 U248 ( .A0(n195), .B0(n194), .CI(\mul_b2/fa1_s2_r[29] ), .CO(
        n393), .S0(n392) );
  HS65_GS_IVX2 U249 ( .A(n392), .Z(n391) );
  HS65_GS_OAI21X2 U250 ( .A(n196), .B(n387), .C(n392), .Z(n821) );
  HS65_GS_PAO2X4 U251 ( .A(\mul_b2/fa1_s1_r[25] ), .B(\mul_b2/fa1_s0_r[25] ), 
        .P(\mul_b2/fa1_c0_r[24] ), .Z(n197) );
  HS65_GSS_XOR2X3 U252 ( .A(n197), .B(\mul_b2/fa1_s2_r[26] ), .Z(n204) );
  HS65_GSS_XOR3X2 U253 ( .A(\mul_b2/fa1_c0_r[25] ), .B(\mul_b2/fa1_s1_r[26] ), 
        .C(\mul_b2/fa1_s0_r[26] ), .Z(n203) );
  HS65_GS_NAND2X2 U254 ( .A(n204), .B(n203), .Z(n202) );
  HS65_GS_IVX2 U255 ( .A(n202), .Z(n199) );
  HS65_GS_AND2X4 U256 ( .A(n197), .B(\mul_b2/fa1_s2_r[26] ), .Z(n198) );
  HS65_GS_OR2X4 U257 ( .A(n199), .B(n198), .Z(n376) );
  HS65_GS_PAO2X4 U258 ( .A(\mul_b2/fa1_c0_r[25] ), .B(\mul_b2/fa1_s1_r[26] ), 
        .P(\mul_b2/fa1_s0_r[26] ), .Z(n377) );
  HS65_GSS_XOR2X3 U259 ( .A(n377), .B(\mul_b2/fa1_s2_r[27] ), .Z(n378) );
  HS65_GSS_XOR3X2 U260 ( .A(\mul_b2/fa1_s1_r[27] ), .B(\mul_b2/fa1_s0_r[27] ), 
        .C(\mul_b2/fa1_c0_r[26] ), .Z(n379) );
  HS65_GS_NAND2X2 U261 ( .A(n378), .B(n379), .Z(n383) );
  HS65_GS_OAI21X2 U262 ( .A(n378), .B(n379), .C(n383), .Z(n375) );
  HS65_GS_NAND2X2 U263 ( .A(n376), .B(n375), .Z(n374) );
  HS65_GS_OAI21X2 U264 ( .A(n199), .B(n198), .C(n374), .Z(n1536) );
  HS65_GSS_XOR3X2 U265 ( .A(\mul_b2/fa1_s1_r[25] ), .B(\mul_b2/fa1_s0_r[25] ), 
        .C(\mul_b2/fa1_c0_r[24] ), .Z(n215) );
  HS65_GS_PAO2X4 U266 ( .A(\mul_b2/fa1_s1_r[24] ), .B(\mul_b2/fa1_s0_r[24] ), 
        .P(\mul_b2/fa1_c0_r[23] ), .Z(n200) );
  HS65_GSS_XOR2X3 U267 ( .A(n200), .B(\mul_b2/fa1_s2_r[25] ), .Z(n216) );
  HS65_GS_AND2X4 U268 ( .A(n200), .B(\mul_b2/fa1_s2_r[25] ), .Z(n201) );
  HS65_GS_AOI12X2 U269 ( .A(n215), .B(n216), .C(n201), .Z(n371) );
  HS65_GS_OAI21X2 U270 ( .A(n204), .B(n203), .C(n202), .Z(n372) );
  HS65_GS_OR2X4 U271 ( .A(n371), .B(n372), .Z(n1789) );
  HS65_GS_PAO2X4 U272 ( .A(\mul_b2/fa1_s1_r[22] ), .B(\mul_b2/fa1_s0_r[22] ), 
        .P(\mul_b2/fa1_c0_r[21] ), .Z(n205) );
  HS65_GSS_XOR3X2 U273 ( .A(\mul_b2/fa1_c0_r[22] ), .B(\mul_b2/fa1_s1_r[23] ), 
        .C(\mul_b2/fa1_s0_r[23] ), .Z(n223) );
  HS65_GS_NAND2X2 U274 ( .A(n224), .B(n223), .Z(n222) );
  HS65_GS_IVX2 U275 ( .A(n222), .Z(n207) );
  HS65_GS_FA1X4 U276 ( .A0(\mul_b2/fa1_s2_r[23] ), .B0(\mul_b2/fa1_c1_r[22] ), 
        .CI(n205), .CO(n206), .S0(n224) );
  HS65_GS_AOI12X2 U277 ( .A(n223), .B(n224), .C(n206), .Z(n208) );
  HS65_GS_AOI13X2 U278 ( .A(n207), .B(\mul_b2/fa1_s2_r[23] ), .C(
        \mul_b2/fa1_c1_r[22] ), .D(n208), .Z(n367) );
  HS65_GS_PAO2X4 U279 ( .A(\mul_b2/fa1_c0_r[22] ), .B(\mul_b2/fa1_s1_r[23] ), 
        .P(\mul_b2/fa1_s0_r[23] ), .Z(n210) );
  HS65_GSS_XOR3X2 U280 ( .A(\mul_b2/fa1_s1_r[24] ), .B(\mul_b2/fa1_s0_r[24] ), 
        .C(\mul_b2/fa1_c0_r[23] ), .Z(n212) );
  HS65_GS_NAND2X2 U281 ( .A(n211), .B(n212), .Z(n209) );
  HS65_GS_OAI21X2 U282 ( .A(n211), .B(n212), .C(n209), .Z(n366) );
  HS65_GS_NAND2X2 U283 ( .A(n367), .B(n366), .Z(n365) );
  HS65_GS_NOR2AX3 U284 ( .A(n365), .B(n208), .Z(n1540) );
  HS65_GS_IVX2 U285 ( .A(n209), .Z(n370) );
  HS65_GS_FA1X4 U286 ( .A0(\mul_b2/fa1_s2_r[24] ), .B0(\mul_b2/fa1_c1_r[23] ), 
        .CI(n210), .CO(n369), .S0(n211) );
  HS65_GS_AOI12X2 U287 ( .A(n212), .B(n211), .C(n369), .Z(n213) );
  HS65_GS_AOI13X2 U288 ( .A(n370), .B(\mul_b2/fa1_c1_r[23] ), .C(
        \mul_b2/fa1_s2_r[24] ), .D(n213), .Z(n218) );
  HS65_GS_NAND2X2 U289 ( .A(n216), .B(n215), .Z(n214) );
  HS65_GS_OAI21X2 U290 ( .A(n216), .B(n215), .C(n214), .Z(n217) );
  HS65_GS_NAND2X2 U291 ( .A(n218), .B(n217), .Z(n368) );
  HS65_GS_OAI21X2 U292 ( .A(n218), .B(n217), .C(n368), .Z(n1539) );
  HS65_GS_PAO2X4 U293 ( .A(\mul_b2/fa1_s1_r[21] ), .B(\mul_b2/fa1_s0_r[21] ), 
        .P(\mul_b2/fa1_c0_r[20] ), .Z(n219) );
  HS65_GSS_XOR3X2 U294 ( .A(\mul_b2/fa1_s1_r[22] ), .B(\mul_b2/fa1_s0_r[22] ), 
        .C(\mul_b2/fa1_c0_r[21] ), .Z(n230) );
  HS65_GS_NAND2X2 U295 ( .A(n231), .B(n230), .Z(n229) );
  HS65_GS_IVX2 U296 ( .A(n229), .Z(n221) );
  HS65_GS_FA1X4 U297 ( .A0(\mul_b2/fa1_s2_r[22] ), .B0(\mul_b2/fa1_c1_r[21] ), 
        .CI(n219), .CO(n220), .S0(n231) );
  HS65_GS_AOI12X2 U298 ( .A(n230), .B(n231), .C(n220), .Z(n225) );
  HS65_GS_AOI13X2 U299 ( .A(n221), .B(\mul_b2/fa1_s2_r[22] ), .C(
        \mul_b2/fa1_c1_r[21] ), .D(n225), .Z(n235) );
  HS65_GS_OAI21X2 U300 ( .A(n224), .B(n223), .C(n222), .Z(n234) );
  HS65_GS_NAND2X2 U301 ( .A(n235), .B(n234), .Z(n233) );
  HS65_GS_NOR2AX3 U302 ( .A(n233), .B(n225), .Z(n1544) );
  HS65_GS_PAO2X4 U303 ( .A(\mul_b2/fa1_s1_r[20] ), .B(\mul_b2/fa1_s0_r[20] ), 
        .P(\mul_b2/fa1_c0_r[19] ), .Z(n226) );
  HS65_GSS_XOR3X2 U304 ( .A(\mul_b2/fa1_s1_r[21] ), .B(\mul_b2/fa1_s0_r[21] ), 
        .C(\mul_b2/fa1_c0_r[20] ), .Z(n240) );
  HS65_GS_NAND2X2 U305 ( .A(n241), .B(n240), .Z(n239) );
  HS65_GS_IVX2 U306 ( .A(n239), .Z(n228) );
  HS65_GS_FA1X4 U307 ( .A0(\mul_b2/fa1_s2_r[21] ), .B0(\mul_b2/fa1_c1_r[20] ), 
        .CI(n226), .CO(n227), .S0(n241) );
  HS65_GS_NOR2X2 U308 ( .A(n228), .B(n227), .Z(n232) );
  HS65_GS_AOI13X2 U309 ( .A(n228), .B(\mul_b2/fa1_s2_r[21] ), .C(
        \mul_b2/fa1_c1_r[20] ), .D(n232), .Z(n364) );
  HS65_GS_OAI21X2 U310 ( .A(n231), .B(n230), .C(n229), .Z(n363) );
  HS65_GS_NAND2X2 U311 ( .A(n364), .B(n363), .Z(n362) );
  HS65_GS_NOR2AX3 U312 ( .A(n362), .B(n232), .Z(n1548) );
  HS65_GS_OAI21X2 U313 ( .A(n235), .B(n234), .C(n233), .Z(n1547) );
  HS65_GS_PAO2X4 U314 ( .A(\mul_b2/fa1_s1_r[19] ), .B(\mul_b2/fa1_s0_r[19] ), 
        .P(\mul_b2/fa1_c0_r[18] ), .Z(n236) );
  HS65_GSS_XOR3X2 U315 ( .A(\mul_b2/fa1_s1_r[20] ), .B(\mul_b2/fa1_s0_r[20] ), 
        .C(\mul_b2/fa1_c0_r[19] ), .Z(n248) );
  HS65_GS_NAND2X2 U316 ( .A(n249), .B(n248), .Z(n247) );
  HS65_GS_IVX2 U317 ( .A(n247), .Z(n238) );
  HS65_GS_FA1X4 U318 ( .A0(\mul_b2/fa1_s2_r[20] ), .B0(\mul_b2/fa1_c1_r[19] ), 
        .CI(n236), .CO(n237), .S0(n249) );
  HS65_GS_AOI12X2 U319 ( .A(n248), .B(n249), .C(n237), .Z(n242) );
  HS65_GS_AOI13X2 U320 ( .A(n238), .B(\mul_b2/fa1_c1_r[19] ), .C(
        \mul_b2/fa1_s2_r[20] ), .D(n242), .Z(n244) );
  HS65_GS_OAI21X2 U321 ( .A(n241), .B(n240), .C(n239), .Z(n243) );
  HS65_GS_AOI12X2 U322 ( .A(n244), .B(n243), .C(n242), .Z(n1552) );
  HS65_GSS_XOR2X3 U323 ( .A(n244), .B(n243), .Z(n843) );
  HS65_GSS_XOR3X2 U324 ( .A(\mul_b2/fa1_s1_r[19] ), .B(\mul_b2/fa1_s0_r[19] ), 
        .C(\mul_b2/fa1_c0_r[18] ), .Z(n257) );
  HS65_GS_NAND2X2 U325 ( .A(n258), .B(n257), .Z(n256) );
  HS65_GS_IVX2 U326 ( .A(n256), .Z(n252) );
  HS65_GS_FA1X4 U327 ( .A0(\mul_b2/fa1_s2_r[19] ), .B0(\mul_b2/fa1_c1_r[18] ), 
        .CI(n245), .CO(n251), .S0(n258) );
  HS65_GS_AOI12X2 U328 ( .A(n257), .B(n258), .C(n251), .Z(n246) );
  HS65_GS_AOI13X2 U329 ( .A(n252), .B(\mul_b2/fa1_c1_r[18] ), .C(
        \mul_b2/fa1_s2_r[19] ), .D(n246), .Z(n361) );
  HS65_GS_OAI21X2 U330 ( .A(n249), .B(n248), .C(n247), .Z(n360) );
  HS65_GS_NAND2X2 U331 ( .A(n361), .B(n360), .Z(n250) );
  HS65_GS_OAI21X2 U332 ( .A(n252), .B(n251), .C(n250), .Z(n841) );
  HS65_GS_FA1X4 U333 ( .A0(\mul_b2/fa1_s0_r[18] ), .B0(\mul_b2/fa1_s1_r[18] ), 
        .CI(\mul_b2/fa1_c0_r[17] ), .CO(n245), .S0(n272) );
  HS65_GS_FA1X4 U334 ( .A0(\mul_b2/fa1_s2_r[18] ), .B0(\mul_b2/fa1_c1_r[17] ), 
        .CI(n253), .CO(n254), .S0(n273) );
  HS65_GS_AOI12X2 U335 ( .A(n272), .B(n273), .C(n254), .Z(n260) );
  HS65_GS_NAND2X2 U336 ( .A(n273), .B(n272), .Z(n271) );
  HS65_GS_IVX2 U337 ( .A(n271), .Z(n255) );
  HS65_GS_AOI13X2 U338 ( .A(n255), .B(\mul_b2/fa1_c1_r[17] ), .C(
        \mul_b2/fa1_s2_r[18] ), .D(n260), .Z(n358) );
  HS65_GS_OAI21X2 U339 ( .A(n258), .B(n257), .C(n256), .Z(n357) );
  HS65_GS_AND2X4 U340 ( .A(n358), .B(n357), .Z(n259) );
  HS65_GS_NOR2X2 U341 ( .A(n260), .B(n259), .Z(n1555) );
  HS65_GS_NAND2X2 U342 ( .A(n280), .B(n279), .Z(n278) );
  HS65_GS_IVX2 U343 ( .A(n278), .Z(n263) );
  HS65_GS_FA1X4 U344 ( .A0(\mul_b2/fa1_s2_r[16] ), .B0(\mul_b2/fa1_c1_r[15] ), 
        .CI(n261), .CO(n262), .S0(n280) );
  HS65_GS_NOR2X2 U345 ( .A(n263), .B(n262), .Z(n264) );
  HS65_GS_AOI13X2 U346 ( .A(n263), .B(\mul_b2/fa1_s2_r[16] ), .C(
        \mul_b2/fa1_c1_r[15] ), .D(n264), .Z(n352) );
  HS65_GS_FA1X4 U347 ( .A0(\mul_b2/fa1_s0_r[16] ), .B0(\mul_b2/fa1_s1_r[16] ), 
        .CI(\mul_b2/fa1_c0_r[15] ), .CO(n266), .S0(n279) );
  HS65_GS_FA1X4 U348 ( .A0(\mul_b2/fa1_s0_r[17] ), .B0(\mul_b2/fa1_s1_r[17] ), 
        .CI(\mul_b2/fa1_c0_r[16] ), .CO(n253), .S0(n269) );
  HS65_GS_NAND2X2 U349 ( .A(n268), .B(n269), .Z(n265) );
  HS65_GS_OAI21X2 U350 ( .A(n268), .B(n269), .C(n265), .Z(n351) );
  HS65_GS_NAND2X2 U351 ( .A(n352), .B(n351), .Z(n350) );
  HS65_GS_NOR2AX3 U352 ( .A(n350), .B(n264), .Z(n1565) );
  HS65_GS_IVX2 U353 ( .A(n265), .Z(n270) );
  HS65_GS_FA1X4 U354 ( .A0(\mul_b2/fa1_s2_r[17] ), .B0(\mul_b2/fa1_c1_r[16] ), 
        .CI(n266), .CO(n267), .S0(n268) );
  HS65_GS_AOI12X2 U355 ( .A(n269), .B(n268), .C(n267), .Z(n353) );
  HS65_GS_AOI13X2 U356 ( .A(n270), .B(\mul_b2/fa1_c1_r[16] ), .C(
        \mul_b2/fa1_s2_r[17] ), .D(n353), .Z(n275) );
  HS65_GS_OAI21X2 U357 ( .A(n273), .B(n272), .C(n271), .Z(n274) );
  HS65_GS_NAND2X2 U358 ( .A(n275), .B(n274), .Z(n354) );
  HS65_GS_OAI21X2 U359 ( .A(n275), .B(n274), .C(n354), .Z(n1564) );
  HS65_GS_AND2X4 U360 ( .A(\mul_b2/fa1_c1_r[14] ), .B(\mul_b2/fa1_s2_r[15] ), 
        .Z(n277) );
  HS65_GS_FA1X4 U361 ( .A0(\mul_b2/fa1_s0_r[15] ), .B0(\mul_b2/fa1_s1_r[15] ), 
        .CI(\mul_b2/fa1_c0_r[14] ), .CO(n261), .S0(n282) );
  HS65_GSS_XOR2X3 U362 ( .A(\mul_b2/fa1_c1_r[14] ), .B(\mul_b2/fa1_s2_r[15] ), 
        .Z(n281) );
  HS65_GS_AOI12X2 U363 ( .A(\mul_b2/fa1_s2_r[15] ), .B(\mul_b2/fa1_c1_r[14] ), 
        .C(n276), .Z(n347) );
  HS65_GS_AOI13X2 U364 ( .A(n277), .B(n282), .C(n283), .D(n347), .Z(n349) );
  HS65_GS_OAI21X2 U365 ( .A(n280), .B(n279), .C(n278), .Z(n348) );
  HS65_GSS_XOR2X3 U366 ( .A(n349), .B(n348), .Z(n846) );
  HS65_GS_FA1X4 U367 ( .A0(n283), .B0(n282), .CI(n281), .CO(n276), .S0(n286)
         );
  HS65_GS_AND2X4 U368 ( .A(\mul_b2/fa1_c1_r[13] ), .B(\mul_b2/fa1_s2_r[14] ), 
        .Z(n285) );
  HS65_GSS_XOR2X3 U369 ( .A(\mul_b2/fa1_c1_r[13] ), .B(\mul_b2/fa1_s2_r[14] ), 
        .Z(n331) );
  HS65_GS_FA1X4 U370 ( .A0(\mul_b2/fa1_s0_r[14] ), .B0(\mul_b2/fa1_s1_r[14] ), 
        .CI(\mul_b2/fa1_c0_r[13] ), .CO(n283), .S0(n330) );
  HS65_GS_FA1X4 U371 ( .A0(n286), .B0(n285), .CI(n284), .CO(n345), .S0(n342)
         );
  HS65_GS_NAND2X2 U372 ( .A(n319), .B(n318), .Z(n317) );
  HS65_GS_IVX2 U373 ( .A(n317), .Z(n289) );
  HS65_GS_FA1X4 U374 ( .A0(\mul_b2/fa1_s2_r[12] ), .B0(\mul_b2/fa1_c1_r[11] ), 
        .CI(n287), .CO(n288), .S0(n319) );
  HS65_GS_AOI12X2 U375 ( .A(n318), .B(n319), .C(n288), .Z(n328) );
  HS65_GS_AOI13X2 U376 ( .A(n289), .B(\mul_b2/fa1_c1_r[11] ), .C(
        \mul_b2/fa1_s2_r[12] ), .D(n328), .Z(n326) );
  HS65_GS_FA1X4 U377 ( .A0(\mul_b2/fa1_s0_r[12] ), .B0(\mul_b2/fa1_s1_r[12] ), 
        .CI(\mul_b2/fa1_c0_r[11] ), .CO(n334), .S0(n318) );
  HS65_GS_FA1X4 U378 ( .A0(\mul_b2/fa1_s0_r[13] ), .B0(\mul_b2/fa1_s1_r[13] ), 
        .CI(\mul_b2/fa1_c0_r[12] ), .CO(n329), .S0(n333) );
  HS65_GSS_XOR2X3 U379 ( .A(\mul_b2/fa1_c1_r[12] ), .B(\mul_b2/fa1_s2_r[13] ), 
        .Z(n332) );
  HS65_GS_FA1X4 U380 ( .A0(\mul_b2/fa1_s0_r[11] ), .B0(\mul_b2/fa1_s1_r[11] ), 
        .CI(\mul_b2/fa1_c0_r[10] ), .CO(n287), .S0(n314) );
  HS65_GS_FA1X4 U381 ( .A0(\mul_b2/fa1_s0_r[10] ), .B0(\mul_b2/fa1_s1_r[10] ), 
        .CI(\mul_b2/fa1_c0_r[9] ), .CO(n315), .S0(n305) );
  HS65_GS_FA1X4 U382 ( .A0(\mul_b2/fa1_s0_r[9] ), .B0(\mul_b2/fa1_s1_r[9] ), 
        .CI(\mul_b2/fa1_c0_r[8] ), .CO(n306), .S0(n310) );
  HS65_GS_PAO2X4 U383 ( .A(\mul_b2/fa1_s1_r[8] ), .B(\mul_b2/fa1_s0_r[8] ), 
        .P(\mul_b2/fa1_c0_r[7] ), .Z(n309) );
  HS65_GS_NOR2X2 U384 ( .A(n309), .B(n310), .Z(n304) );
  HS65_GSS_XOR3X2 U385 ( .A(\mul_b2/fa1_s1_r[8] ), .B(\mul_b2/fa1_s0_r[8] ), 
        .C(\mul_b2/fa1_c0_r[7] ), .Z(n302) );
  HS65_GS_PAO2X4 U386 ( .A(\mul_b2/fa1_c0_r[6] ), .B(\mul_b2/fa1_s1_r[7] ), 
        .P(\mul_b2/fa1_s0_r[7] ), .Z(n301) );
  HS65_GS_PAO2X4 U387 ( .A(\mul_b2/fa1_s1_r[6] ), .B(\mul_b2/fa1_s0_r[6] ), 
        .P(\mul_b2/fa1_c0_r[5] ), .Z(n299) );
  HS65_GSS_XOR3X2 U388 ( .A(\mul_b2/fa1_c0_r[6] ), .B(\mul_b2/fa1_s1_r[7] ), 
        .C(\mul_b2/fa1_s0_r[7] ), .Z(n298) );
  HS65_GS_NOR2X2 U389 ( .A(n299), .B(n298), .Z(n296) );
  HS65_GS_AND2X4 U390 ( .A(\mul_b2/fa1_c0_r[4] ), .B(\mul_b2/fa1_s0_r[5] ), 
        .Z(n294) );
  HS65_GSS_XOR3X2 U391 ( .A(\mul_b2/fa1_s1_r[6] ), .B(\mul_b2/fa1_s0_r[6] ), 
        .C(\mul_b2/fa1_c0_r[5] ), .Z(n293) );
  HS65_GSS_XOR2X3 U392 ( .A(\mul_b2/fa1_c0_r[4] ), .B(\mul_b2/fa1_s0_r[5] ), 
        .Z(n291) );
  HS65_GS_AND2X4 U393 ( .A(\mul_b2/fa1_c0_r[3] ), .B(\mul_b2/fa1_s0_r[4] ), 
        .Z(n290) );
  HS65_GS_AND2X4 U394 ( .A(n291), .B(n290), .Z(n292) );
  HS65_GS_PAOI2X1 U395 ( .A(n294), .B(n293), .P(n292), .Z(n295) );
  HS65_GS_NOR2X2 U396 ( .A(n296), .B(n295), .Z(n297) );
  HS65_GS_AO12X4 U397 ( .A(n299), .B(n298), .C(n297), .Z(n300) );
  HS65_GS_PAOI2X1 U398 ( .A(n302), .B(n301), .P(n300), .Z(n303) );
  HS65_GS_NOR2X2 U399 ( .A(n304), .B(n303), .Z(n308) );
  HS65_GS_FA1X4 U400 ( .A0(\mul_b2/fa1_c1_r[9] ), .B0(n306), .CI(n305), .CO(
        n312), .S0(n307) );
  HS65_GS_CB4I1X4 U401 ( .A(n310), .B(n309), .C(n308), .D(n307), .Z(n311) );
  HS65_GS_PAOI2X1 U402 ( .A(n313), .B(n312), .P(n311), .Z(n322) );
  HS65_GS_FA1X4 U403 ( .A0(\mul_b2/fa1_c1_r[10] ), .B0(n315), .CI(n314), .CO(
        n316), .S0(n313) );
  HS65_GS_IVX2 U404 ( .A(n316), .Z(n321) );
  HS65_GS_OAI21X2 U405 ( .A(n319), .B(n318), .C(n317), .Z(n320) );
  HS65_GS_PAOI2X1 U406 ( .A(n322), .B(n321), .P(n320), .Z(n323) );
  HS65_GS_OAI21X2 U407 ( .A(n326), .B(n325), .C(n323), .Z(n324) );
  HS65_GS_AOI12X2 U408 ( .A(n326), .B(n325), .C(n324), .Z(n336) );
  HS65_GS_NOR2AX3 U409 ( .A(n326), .B(n325), .Z(n327) );
  HS65_GS_NOR2X2 U410 ( .A(n328), .B(n327), .Z(n335) );
  HS65_GS_NAND2X2 U411 ( .A(n336), .B(n335), .Z(n337) );
  HS65_GS_AND2X4 U412 ( .A(\mul_b2/fa1_c1_r[12] ), .B(\mul_b2/fa1_s2_r[13] ), 
        .Z(n340) );
  HS65_GS_FA1X4 U413 ( .A0(n331), .B0(n330), .CI(n329), .CO(n284), .S0(n339)
         );
  HS65_GS_FA1X4 U414 ( .A0(n334), .B0(n333), .CI(n332), .CO(n338), .S0(n325)
         );
  HS65_GSS_XOR2X3 U415 ( .A(n336), .B(n335), .Z(n1578) );
  HS65_GS_NAND2X2 U416 ( .A(n1579), .B(n1578), .Z(n1577) );
  HS65_GS_NAND2X2 U417 ( .A(n337), .B(n1577), .Z(n341) );
  HS65_GS_NAND2X2 U418 ( .A(n342), .B(n341), .Z(n343) );
  HS65_GS_FA1X4 U419 ( .A0(n340), .B0(n339), .CI(n338), .CO(n1575), .S0(n1579)
         );
  HS65_GSS_XOR2X3 U420 ( .A(n342), .B(n341), .Z(n1574) );
  HS65_GS_NAND2X2 U421 ( .A(n1575), .B(n1574), .Z(n1573) );
  HS65_GS_NAND2X2 U422 ( .A(n343), .B(n1573), .Z(n344) );
  HS65_GSS_XNOR2X3 U423 ( .A(n345), .B(n344), .Z(n847) );
  HS65_GS_NAND2X2 U424 ( .A(n345), .B(n344), .Z(n346) );
  HS65_GS_OAI21X2 U425 ( .A(n846), .B(n847), .C(n346), .Z(n1569) );
  HS65_GS_AOI12X2 U426 ( .A(n349), .B(n348), .C(n347), .Z(n1568) );
  HS65_GS_OAI21X2 U427 ( .A(n352), .B(n351), .C(n350), .Z(n1567) );
  HS65_GS_NOR2AX3 U428 ( .A(n354), .B(n353), .Z(n355) );
  HS65_GS_NAND2X2 U429 ( .A(n356), .B(n355), .Z(n359) );
  HS65_GSS_XOR2X3 U430 ( .A(n356), .B(n355), .Z(n1561) );
  HS65_GSS_XNOR2X3 U431 ( .A(n358), .B(n357), .Z(n1560) );
  HS65_GS_NAND2X2 U432 ( .A(n1561), .B(n1560), .Z(n1559) );
  HS65_GS_NAND2X2 U433 ( .A(n359), .B(n1559), .Z(n1554) );
  HS65_GSS_XNOR2X3 U434 ( .A(n361), .B(n360), .Z(n1557) );
  HS65_GS_PAOI2X1 U435 ( .A(n1555), .B(n1554), .P(n1557), .Z(n840) );
  HS65_GS_PAOI2X1 U436 ( .A(n843), .B(n841), .P(n840), .Z(n1551) );
  HS65_GS_OAI21X2 U437 ( .A(n364), .B(n363), .C(n362), .Z(n1550) );
  HS65_GS_OAI21X2 U438 ( .A(n367), .B(n366), .C(n365), .Z(n1542) );
  HS65_GS_OA12X4 U439 ( .A(n370), .B(n369), .C(n368), .Z(n816) );
  HS65_GS_IVX2 U440 ( .A(n371), .Z(n373) );
  HS65_GSS_XNOR2X3 U441 ( .A(n373), .B(n372), .Z(n818) );
  HS65_GS_PAOI2X1 U442 ( .A(n817), .B(n816), .P(n818), .Z(n1788) );
  HS65_GS_OA12X4 U443 ( .A(n376), .B(n375), .C(n374), .Z(n1787) );
  HS65_GS_AND2X4 U444 ( .A(\mul_b2/fa1_s2_r[27] ), .B(n377), .Z(n385) );
  HS65_GS_AO12X4 U445 ( .A(n379), .B(n378), .C(n385), .Z(n382) );
  HS65_GS_OAI21X2 U446 ( .A(n388), .B(n389), .C(n380), .Z(n381) );
  HS65_GS_NAND2X2 U447 ( .A(n382), .B(n381), .Z(n384) );
  HS65_GS_OA12X4 U448 ( .A(n382), .B(n381), .C(n384), .Z(n1534) );
  HS65_GS_IVX2 U449 ( .A(n383), .Z(n386) );
  HS65_GS_OAI21X2 U450 ( .A(n386), .B(n385), .C(n384), .Z(n826) );
  HS65_GS_AO12X4 U451 ( .A(n389), .B(n388), .C(n387), .Z(n390) );
  HS65_GS_MUXI21X2 U452 ( .D0(n392), .D1(n391), .S0(n390), .Z(n825) );
  HS65_GS_MUXI21X2 U453 ( .D0(n395), .D1(n394), .S0(n393), .Z(n819) );
  HS65_GS_FA1X4 U454 ( .A0(n397), .B0(n396), .CI(\mul_b2/fa1_s2_r[30] ), .CO(
        n400), .S0(n395) );
  HS65_GS_FA1X4 U455 ( .A0(\mul_b2/fa1_s2_r[31] ), .B0(n399), .CI(n398), .CO(
        n192), .S0(n401) );
  HS65_GSS_XNOR2X3 U456 ( .A(n400), .B(n401), .Z(n822) );
  HS65_GS_NAND2X2 U457 ( .A(n401), .B(n400), .Z(n828) );
  HS65_GSS_XOR2X3 U458 ( .A(n403), .B(n402), .Z(n404) );
  HS65_GSS_XOR2X3 U459 ( .A(n405), .B(n404), .Z(n406) );
  HS65_GSS_XNOR2X3 U460 ( .A(n406), .B(\mul_b2/fa1_c0_r[32] ), .Z(n407) );
  HS65_GSS_XOR3X2 U461 ( .A(n407), .B(\mul_b2/fa1_s0_r[33] ), .C(
        \mul_b2/fa1_s1_r[33] ), .Z(n408) );
  HS65_GSS_XOR3X2 U462 ( .A(n409), .B(\mul_b2/fa1_s2_r[33] ), .C(n408), .Z(
        \mul_b2/result_sat[15] ) );
  HS65_GS_IVX2 U463 ( .A(x_z2[15]), .Z(n1439) );
  HS65_GS_IVX4 U464 ( .A(n1439), .Z(\DP_OP_331J1_157_5454/n87 ) );
  HS65_GS_IVX2 U465 ( .A(y_z1[15]), .Z(n1705) );
  HS65_GS_IVX2 U466 ( .A(x_reg2[15]), .Z(n1494) );
  HS65_GS_IVX4 U467 ( .A(n1494), .Z(\DP_OP_371J1_181_1383/n79 ) );
  HS65_GS_PAO2X4 U468 ( .A(\mul_b1/fa1_c0_r[31] ), .B(\mul_b1/fa1_s1_r[32] ), 
        .P(\mul_b1/fa1_s0_r[32] ), .Z(n614) );
  HS65_GS_AND2X4 U469 ( .A(\mul_b1/fa1_c1_r[31] ), .B(\mul_b1/fa1_s2_r[32] ), 
        .Z(n613) );
  HS65_GSS_XOR2X3 U470 ( .A(\mul_b1/fa1_s2_r[32] ), .B(\mul_b1/fa1_c1_r[31] ), 
        .Z(n412) );
  HS65_GSS_XOR3X2 U471 ( .A(\mul_b1/fa1_c0_r[31] ), .B(\mul_b1/fa1_s1_r[32] ), 
        .C(\mul_b1/fa1_s0_r[32] ), .Z(n411) );
  HS65_GS_PAO2X4 U472 ( .A(\mul_b1/fa1_c0_r[30] ), .B(\mul_b1/fa1_s1_r[31] ), 
        .P(\mul_b1/fa1_s0_r[31] ), .Z(n410) );
  HS65_GS_AND2X4 U473 ( .A(\mul_b1/fa1_s2_r[31] ), .B(\mul_b1/fa1_c1_r[30] ), 
        .Z(n415) );
  HS65_GSS_XOR2X3 U474 ( .A(\mul_b1/fa1_s2_r[31] ), .B(\mul_b1/fa1_c1_r[30] ), 
        .Z(n602) );
  HS65_GSS_XOR3X2 U475 ( .A(\mul_b1/fa1_c0_r[30] ), .B(\mul_b1/fa1_s1_r[31] ), 
        .C(\mul_b1/fa1_s0_r[31] ), .Z(n601) );
  HS65_GS_PAO2X4 U476 ( .A(\mul_b1/fa1_c0_r[29] ), .B(\mul_b1/fa1_s1_r[30] ), 
        .P(\mul_b1/fa1_s0_r[30] ), .Z(n600) );
  HS65_GS_FA1X4 U477 ( .A0(n412), .B0(n411), .CI(n410), .CO(n611), .S0(n413)
         );
  HS65_GS_FA1X4 U478 ( .A0(n415), .B0(n414), .CI(n413), .CO(n610), .S0(n1039)
         );
  HS65_GS_FA1X4 U479 ( .A0(\mul_b1/fa1_c1_r[27] ), .B0(\mul_b1/fa1_c2_r[27] ), 
        .CI(\mul_b1/fa1_s2_r[28] ), .CO(n590), .S0(n584) );
  HS65_GS_PAO2X4 U480 ( .A(\mul_b1/fa1_c0_r[26] ), .B(\mul_b1/fa1_s1_r[27] ), 
        .P(\mul_b1/fa1_s0_r[27] ), .Z(n583) );
  HS65_GSS_XOR3X2 U481 ( .A(\mul_b1/fa1_c0_r[27] ), .B(\mul_b1/fa1_s1_r[28] ), 
        .C(\mul_b1/fa1_s0_r[28] ), .Z(n582) );
  HS65_GS_PAO2X4 U482 ( .A(\mul_b1/fa1_c0_r[27] ), .B(\mul_b1/fa1_s1_r[28] ), 
        .P(\mul_b1/fa1_s0_r[28] ), .Z(n592) );
  HS65_GSS_XOR3X2 U483 ( .A(\mul_b1/fa1_c0_r[28] ), .B(\mul_b1/fa1_s1_r[29] ), 
        .C(\mul_b1/fa1_s0_r[29] ), .Z(n591) );
  HS65_GS_FA1X4 U484 ( .A0(\mul_b1/fa1_c1_r[25] ), .B0(\mul_b1/fa1_c2_r[25] ), 
        .CI(\mul_b1/fa1_s2_r[26] ), .CO(n578), .S0(n418) );
  HS65_GS_PAO2X4 U485 ( .A(\mul_b1/fa1_s1_r[25] ), .B(\mul_b1/fa1_s0_r[25] ), 
        .P(\mul_b1/fa1_c0_r[24] ), .Z(n417) );
  HS65_GSS_XOR3X2 U486 ( .A(\mul_b1/fa1_c0_r[25] ), .B(\mul_b1/fa1_s1_r[26] ), 
        .C(\mul_b1/fa1_s0_r[26] ), .Z(n416) );
  HS65_GS_PAO2X4 U487 ( .A(\mul_b1/fa1_c0_r[25] ), .B(\mul_b1/fa1_s1_r[26] ), 
        .P(\mul_b1/fa1_s0_r[26] ), .Z(n580) );
  HS65_GSS_XOR3X2 U488 ( .A(\mul_b1/fa1_c0_r[26] ), .B(\mul_b1/fa1_s1_r[27] ), 
        .C(\mul_b1/fa1_s0_r[27] ), .Z(n579) );
  HS65_GS_FA1X4 U489 ( .A0(\mul_b1/fa1_c1_r[24] ), .B0(\mul_b1/fa1_c2_r[24] ), 
        .CI(\mul_b1/fa1_s2_r[25] ), .CO(n575), .S0(n569) );
  HS65_GS_PAO2X4 U490 ( .A(\mul_b1/fa1_c0_r[23] ), .B(\mul_b1/fa1_s1_r[24] ), 
        .P(\mul_b1/fa1_s0_r[24] ), .Z(n568) );
  HS65_GSS_XOR3X2 U491 ( .A(\mul_b1/fa1_s1_r[25] ), .B(\mul_b1/fa1_s0_r[25] ), 
        .C(\mul_b1/fa1_c0_r[24] ), .Z(n567) );
  HS65_GS_FA1X4 U492 ( .A0(n418), .B0(n417), .CI(n416), .CO(n577), .S0(n573)
         );
  HS65_GS_FA1X4 U493 ( .A0(\mul_b1/fa1_c1_r[21] ), .B0(\mul_b1/fa1_c2_r[21] ), 
        .CI(\mul_b1/fa1_s2_r[22] ), .CO(n557), .S0(n421) );
  HS65_GS_PAO2X4 U494 ( .A(\mul_b1/fa1_s1_r[21] ), .B(\mul_b1/fa1_s0_r[21] ), 
        .P(\mul_b1/fa1_c0_r[20] ), .Z(n420) );
  HS65_GSS_XOR3X2 U495 ( .A(\mul_b1/fa1_c0_r[21] ), .B(\mul_b1/fa1_s1_r[22] ), 
        .C(\mul_b1/fa1_s0_r[22] ), .Z(n419) );
  HS65_GS_PAO2X4 U496 ( .A(\mul_b1/fa1_c0_r[21] ), .B(\mul_b1/fa1_s1_r[22] ), 
        .P(\mul_b1/fa1_s0_r[22] ), .Z(n559) );
  HS65_GSS_XOR3X2 U497 ( .A(\mul_b1/fa1_c0_r[22] ), .B(\mul_b1/fa1_s1_r[23] ), 
        .C(\mul_b1/fa1_s0_r[23] ), .Z(n558) );
  HS65_GS_FA1X4 U498 ( .A0(\mul_b1/fa1_c1_r[20] ), .B0(\mul_b1/fa1_c2_r[20] ), 
        .CI(\mul_b1/fa1_s2_r[21] ), .CO(n554), .S0(n548) );
  HS65_GS_PAO2X4 U499 ( .A(\mul_b1/fa1_c0_r[19] ), .B(\mul_b1/fa1_s1_r[20] ), 
        .P(\mul_b1/fa1_s0_r[20] ), .Z(n547) );
  HS65_GSS_XOR3X2 U500 ( .A(\mul_b1/fa1_s1_r[21] ), .B(\mul_b1/fa1_s0_r[21] ), 
        .C(\mul_b1/fa1_c0_r[20] ), .Z(n546) );
  HS65_GS_FA1X4 U501 ( .A0(n421), .B0(n420), .CI(n419), .CO(n556), .S0(n552)
         );
  HS65_GS_FA1X4 U502 ( .A0(\mul_b1/fa1_c1_r[18] ), .B0(\mul_b1/fa1_c2_r[18] ), 
        .CI(\mul_b1/fa1_s2_r[19] ), .CO(n542), .S0(n424) );
  HS65_GS_PAO2X4 U503 ( .A(\mul_b1/fa1_s1_r[18] ), .B(\mul_b1/fa1_s0_r[18] ), 
        .P(\mul_b1/fa1_c0_r[17] ), .Z(n423) );
  HS65_GSS_XOR3X2 U504 ( .A(\mul_b1/fa1_c0_r[18] ), .B(\mul_b1/fa1_s1_r[19] ), 
        .C(\mul_b1/fa1_s0_r[19] ), .Z(n422) );
  HS65_GS_PAO2X4 U505 ( .A(\mul_b1/fa1_c0_r[18] ), .B(\mul_b1/fa1_s1_r[19] ), 
        .P(\mul_b1/fa1_s0_r[19] ), .Z(n544) );
  HS65_GSS_XOR3X2 U506 ( .A(\mul_b1/fa1_c0_r[19] ), .B(\mul_b1/fa1_s1_r[20] ), 
        .C(\mul_b1/fa1_s0_r[20] ), .Z(n543) );
  HS65_GS_FA1X4 U507 ( .A0(\mul_b1/fa1_c1_r[17] ), .B0(\mul_b1/fa1_c2_r[17] ), 
        .CI(\mul_b1/fa1_s2_r[18] ), .CO(n539), .S0(n427) );
  HS65_GS_PAO2X4 U508 ( .A(\mul_b1/fa1_s1_r[17] ), .B(\mul_b1/fa1_s0_r[17] ), 
        .P(\mul_b1/fa1_c0_r[16] ), .Z(n426) );
  HS65_GSS_XOR3X2 U509 ( .A(\mul_b1/fa1_s1_r[18] ), .B(\mul_b1/fa1_s0_r[18] ), 
        .C(\mul_b1/fa1_c0_r[17] ), .Z(n425) );
  HS65_GS_FA1X4 U510 ( .A0(n424), .B0(n423), .CI(n422), .CO(n541), .S0(n537)
         );
  HS65_GS_FA1X4 U511 ( .A0(\mul_b1/fa1_c1_r[16] ), .B0(\mul_b1/fa1_c2_r[16] ), 
        .CI(\mul_b1/fa1_s2_r[17] ), .CO(n536), .S0(n430) );
  HS65_GSS_XOR3X2 U512 ( .A(\mul_b1/fa1_s1_r[17] ), .B(\mul_b1/fa1_s0_r[17] ), 
        .C(\mul_b1/fa1_c0_r[16] ), .Z(n428) );
  HS65_GS_FA1X4 U513 ( .A0(n427), .B0(n426), .CI(n425), .CO(n538), .S0(n534)
         );
  HS65_GS_FA1X4 U514 ( .A0(\mul_b1/fa1_c1_r[15] ), .B0(\mul_b1/fa1_c2_r[15] ), 
        .CI(\mul_b1/fa1_s2_r[16] ), .CO(n533), .S0(n527) );
  HS65_GS_FA1X4 U515 ( .A0(\mul_b1/fa1_s0_r[16] ), .B0(\mul_b1/fa1_s1_r[16] ), 
        .CI(\mul_b1/fa1_c0_r[15] ), .CO(n429), .S0(n525) );
  HS65_GS_FA1X4 U516 ( .A0(n430), .B0(n429), .CI(n428), .CO(n535), .S0(n531)
         );
  HS65_GS_AND2X4 U517 ( .A(\mul_b1/fa1_c1_r[13] ), .B(\mul_b1/fa1_s2_r[14] ), 
        .Z(n521) );
  HS65_GS_FA1X4 U518 ( .A0(\mul_b1/fa1_s0_r[15] ), .B0(\mul_b1/fa1_s1_r[15] ), 
        .CI(\mul_b1/fa1_c0_r[14] ), .CO(n526), .S0(n524) );
  HS65_GSS_XOR2X3 U519 ( .A(\mul_b1/fa1_c1_r[13] ), .B(\mul_b1/fa1_s2_r[14] ), 
        .Z(n510) );
  HS65_GS_FA1X4 U520 ( .A0(\mul_b1/fa1_s0_r[14] ), .B0(\mul_b1/fa1_s1_r[14] ), 
        .CI(\mul_b1/fa1_c0_r[13] ), .CO(n522), .S0(n509) );
  HS65_GS_PAO2X4 U521 ( .A(\mul_b1/fa1_s1_r[11] ), .B(\mul_b1/fa1_c0_r[10] ), 
        .P(\mul_b1/fa1_s0_r[11] ), .Z(n431) );
  HS65_GSS_XOR2X3 U522 ( .A(\mul_b1/fa1_c1_r[11] ), .B(n431), .Z(n439) );
  HS65_GS_NAND2X2 U523 ( .A(n438), .B(n439), .Z(n437) );
  HS65_GS_NAND2X2 U524 ( .A(\mul_b1/fa1_c1_r[11] ), .B(n431), .Z(n432) );
  HS65_GS_NAND2X2 U525 ( .A(n437), .B(n432), .Z(n503) );
  HS65_GS_IVX2 U526 ( .A(n503), .Z(n434) );
  HS65_GS_FA1X4 U527 ( .A0(\mul_b1/fa1_s0_r[13] ), .B0(\mul_b1/fa1_s1_r[13] ), 
        .CI(\mul_b1/fa1_c0_r[12] ), .CO(n508), .S0(n513) );
  HS65_GSS_XOR2X3 U528 ( .A(\mul_b1/fa1_s2_r[13] ), .B(\mul_b1/fa1_c1_r[12] ), 
        .Z(n512) );
  HS65_GS_FA1X4 U529 ( .A0(\mul_b1/fa1_s0_r[12] ), .B0(\mul_b1/fa1_s1_r[12] ), 
        .CI(\mul_b1/fa1_c0_r[11] ), .CO(n511), .S0(n438) );
  HS65_GS_IVX2 U530 ( .A(n433), .Z(n504) );
  HS65_GS_OR2X4 U531 ( .A(n434), .B(n504), .Z(n1795) );
  HS65_GSS_XOR3X2 U532 ( .A(\mul_b1/fa1_s1_r[11] ), .B(\mul_b1/fa1_c0_r[10] ), 
        .C(\mul_b1/fa1_s0_r[11] ), .Z(n489) );
  HS65_GS_PAO2X4 U533 ( .A(\mul_b1/fa1_s0_r[10] ), .B(\mul_b1/fa1_c0_r[9] ), 
        .P(\mul_b1/fa1_s1_r[10] ), .Z(n435) );
  HS65_GSS_XOR2X3 U534 ( .A(\mul_b1/fa1_c1_r[10] ), .B(n435), .Z(n490) );
  HS65_GS_NAND2X2 U535 ( .A(n489), .B(n490), .Z(n488) );
  HS65_GS_NAND2X2 U536 ( .A(\mul_b1/fa1_c1_r[10] ), .B(n435), .Z(n436) );
  HS65_GS_NAND2X2 U537 ( .A(n488), .B(n436), .Z(n442) );
  HS65_GS_IVX2 U538 ( .A(n442), .Z(n440) );
  HS65_GS_OAI21X2 U539 ( .A(n439), .B(n438), .C(n437), .Z(n441) );
  HS65_GS_NOR2X2 U540 ( .A(n440), .B(n441), .Z(n507) );
  HS65_GSS_XOR2X3 U541 ( .A(n442), .B(n441), .Z(n502) );
  HS65_GSS_XOR3X2 U542 ( .A(\mul_b1/fa1_s1_r[9] ), .B(\mul_b1/fa1_c0_r[8] ), 
        .C(\mul_b1/fa1_s0_r[9] ), .Z(n474) );
  HS65_GS_PAO2X4 U543 ( .A(\mul_b1/fa1_s0_r[8] ), .B(\mul_b1/fa1_c0_r[7] ), 
        .P(\mul_b1/fa1_s1_r[8] ), .Z(n443) );
  HS65_GSS_XOR2X3 U544 ( .A(\mul_b1/fa1_c1_r[8] ), .B(n443), .Z(n475) );
  HS65_GS_NAND2X2 U545 ( .A(n474), .B(n475), .Z(n473) );
  HS65_GS_NAND2X2 U546 ( .A(\mul_b1/fa1_c1_r[8] ), .B(n443), .Z(n444) );
  HS65_GS_NAND2X2 U547 ( .A(n473), .B(n444), .Z(n449) );
  HS65_GS_IVX2 U548 ( .A(n449), .Z(n447) );
  HS65_GS_PAOI2X1 U549 ( .A(\mul_b1/fa1_s1_r[9] ), .B(\mul_b1/fa1_c0_r[8] ), 
        .P(\mul_b1/fa1_s0_r[9] ), .Z(n485) );
  HS65_GSS_XNOR2X3 U550 ( .A(\mul_b1/fa1_c1_r[9] ), .B(n485), .Z(n446) );
  HS65_GSS_XOR3X2 U551 ( .A(\mul_b1/fa1_s0_r[10] ), .B(\mul_b1/fa1_c0_r[9] ), 
        .C(\mul_b1/fa1_s1_r[10] ), .Z(n445) );
  HS65_GS_NAND2X2 U552 ( .A(n445), .B(n446), .Z(n495) );
  HS65_GS_OAI21X2 U553 ( .A(n446), .B(n445), .C(n495), .Z(n448) );
  HS65_GS_NOR2X2 U554 ( .A(n447), .B(n448), .Z(n494) );
  HS65_GSS_XOR2X3 U555 ( .A(n449), .B(n448), .Z(n484) );
  HS65_GSS_XOR3X2 U556 ( .A(\mul_b1/fa1_s1_r[7] ), .B(\mul_b1/fa1_c0_r[6] ), 
        .C(\mul_b1/fa1_s0_r[7] ), .Z(n461) );
  HS65_GS_PAO2X4 U557 ( .A(\mul_b1/fa1_s0_r[6] ), .B(\mul_b1/fa1_c0_r[5] ), 
        .P(\mul_b1/fa1_s1_r[6] ), .Z(n462) );
  HS65_GS_NAND2X2 U558 ( .A(n461), .B(n462), .Z(n460) );
  HS65_GS_PAO2X4 U559 ( .A(\mul_b1/fa1_s1_r[7] ), .B(\mul_b1/fa1_c0_r[6] ), 
        .P(\mul_b1/fa1_s0_r[7] ), .Z(n451) );
  HS65_GSS_XOR3X2 U560 ( .A(\mul_b1/fa1_s0_r[8] ), .B(\mul_b1/fa1_c0_r[7] ), 
        .C(\mul_b1/fa1_s1_r[8] ), .Z(n450) );
  HS65_GS_NAND2X2 U561 ( .A(n450), .B(n451), .Z(n479) );
  HS65_GS_OAI21X2 U562 ( .A(n451), .B(n450), .C(n479), .Z(n472) );
  HS65_GS_NOR2X2 U563 ( .A(n460), .B(n472), .Z(n478) );
  HS65_GSS_XOR2X3 U564 ( .A(\mul_b1/fa1_c0_r[4] ), .B(\mul_b1/fa1_s0_r[5] ), 
        .Z(n456) );
  HS65_GS_AND2X4 U565 ( .A(\mul_b1/fa1_s0_r[4] ), .B(\mul_b1/fa1_c0_r[3] ), 
        .Z(n452) );
  HS65_GS_NAND2X2 U566 ( .A(n456), .B(n452), .Z(n453) );
  HS65_GSS_XOR3X2 U567 ( .A(\mul_b1/fa1_s0_r[6] ), .B(\mul_b1/fa1_c0_r[5] ), 
        .C(\mul_b1/fa1_s1_r[6] ), .Z(n467) );
  HS65_GS_IVX2 U568 ( .A(n467), .Z(n459) );
  HS65_GS_NOR2X2 U569 ( .A(n453), .B(n459), .Z(n465) );
  HS65_GS_AND2X4 U570 ( .A(\mul_b1/fa1_c0_r[2] ), .B(\mul_b1/fa1_s0_r[3] ), 
        .Z(n455) );
  HS65_GSS_XOR2X3 U571 ( .A(\mul_b1/fa1_c0_r[3] ), .B(\mul_b1/fa1_s0_r[4] ), 
        .Z(n454) );
  HS65_GS_AND2X4 U572 ( .A(n455), .B(n454), .Z(n457) );
  HS65_GS_NAND2X2 U573 ( .A(n457), .B(n456), .Z(n458) );
  HS65_GS_NOR2X2 U574 ( .A(n459), .B(n458), .Z(n464) );
  HS65_GS_OAI21X2 U575 ( .A(n462), .B(n461), .C(n460), .Z(n463) );
  HS65_GS_IVX2 U576 ( .A(n463), .Z(n468) );
  HS65_GS_PAOI2X1 U577 ( .A(n465), .B(n464), .P(n468), .Z(n471) );
  HS65_GS_AND2X4 U578 ( .A(\mul_b1/fa1_c0_r[4] ), .B(\mul_b1/fa1_s0_r[5] ), 
        .Z(n466) );
  HS65_GS_AND2X4 U579 ( .A(n467), .B(n466), .Z(n469) );
  HS65_GS_NAND2X2 U580 ( .A(n469), .B(n468), .Z(n470) );
  HS65_GS_PAOI2X1 U581 ( .A(n472), .B(n471), .P(n470), .Z(n477) );
  HS65_GS_OAI21X2 U582 ( .A(n475), .B(n474), .C(n473), .Z(n476) );
  HS65_GS_IVX2 U583 ( .A(n476), .Z(n480) );
  HS65_GS_PAOI2X1 U584 ( .A(n478), .B(n477), .P(n480), .Z(n483) );
  HS65_GS_IVX2 U585 ( .A(n479), .Z(n481) );
  HS65_GS_NAND2X2 U586 ( .A(n481), .B(n480), .Z(n482) );
  HS65_GS_PAOI2X1 U587 ( .A(n484), .B(n483), .P(n482), .Z(n493) );
  HS65_GS_IVX2 U588 ( .A(\mul_b1/fa1_c1_r[9] ), .Z(n486) );
  HS65_GS_NOR2X2 U589 ( .A(n486), .B(n485), .Z(n498) );
  HS65_GS_IVX2 U590 ( .A(n498), .Z(n487) );
  HS65_GS_NAND2X2 U591 ( .A(n487), .B(n495), .Z(n491) );
  HS65_GS_OAI21X2 U592 ( .A(n490), .B(n489), .C(n488), .Z(n496) );
  HS65_GSS_XNOR2X3 U593 ( .A(n491), .B(n496), .Z(n492) );
  HS65_GS_PAOI2X1 U594 ( .A(n494), .B(n493), .P(n492), .Z(n501) );
  HS65_GS_IVX2 U595 ( .A(n495), .Z(n499) );
  HS65_GS_IVX2 U596 ( .A(n496), .Z(n497) );
  HS65_GS_OAI21X2 U597 ( .A(n499), .B(n498), .C(n497), .Z(n500) );
  HS65_GS_PAOI2X1 U598 ( .A(n502), .B(n501), .P(n500), .Z(n506) );
  HS65_GSS_XNOR2X3 U599 ( .A(n504), .B(n503), .Z(n505) );
  HS65_GS_PAOI2X1 U600 ( .A(n507), .B(n506), .P(n505), .Z(n1794) );
  HS65_GS_AND2X4 U601 ( .A(\mul_b1/fa1_s2_r[13] ), .B(\mul_b1/fa1_c1_r[12] ), 
        .Z(n518) );
  HS65_GS_FA1X4 U602 ( .A0(n510), .B0(n509), .CI(n508), .CO(n519), .S0(n517)
         );
  HS65_GS_FA1X4 U603 ( .A0(n513), .B0(n512), .CI(n511), .CO(n516), .S0(n433)
         );
  HS65_GS_IVX2 U604 ( .A(n514), .Z(n1793) );
  HS65_GS_IVX2 U605 ( .A(n515), .Z(n1100) );
  HS65_GS_FA1X4 U606 ( .A0(n518), .B0(n517), .CI(n516), .CO(n1099), .S0(n514)
         );
  HS65_GS_FA1X4 U607 ( .A0(n521), .B0(n520), .CI(n519), .CO(n1096), .S0(n1101)
         );
  HS65_GS_FA1X4 U608 ( .A0(\mul_b1/fa1_c1_r[14] ), .B0(\mul_b1/fa1_c2_r[14] ), 
        .CI(\mul_b1/fa1_s2_r[15] ), .CO(n530), .S0(n523) );
  HS65_GS_FA1X4 U609 ( .A0(n524), .B0(n523), .CI(n522), .CO(n529), .S0(n520)
         );
  HS65_GS_FA1X4 U610 ( .A0(n527), .B0(n526), .CI(n525), .CO(n532), .S0(n528)
         );
  HS65_GS_FA1X4 U611 ( .A0(n530), .B0(n529), .CI(n528), .CO(n1092), .S0(n1095)
         );
  HS65_GS_FA1X4 U612 ( .A0(n533), .B0(n532), .CI(n531), .CO(n1089), .S0(n1091)
         );
  HS65_GS_FA1X4 U613 ( .A0(n536), .B0(n535), .CI(n534), .CO(n1085), .S0(n1087)
         );
  HS65_GS_FA1X4 U614 ( .A0(n539), .B0(n538), .CI(n537), .CO(n1081), .S0(n1083)
         );
  HS65_GS_FA1X4 U615 ( .A0(n542), .B0(n541), .CI(n540), .CO(n1077), .S0(n1079)
         );
  HS65_GS_FA1X4 U616 ( .A0(\mul_b1/fa1_c1_r[19] ), .B0(\mul_b1/fa1_c2_r[19] ), 
        .CI(\mul_b1/fa1_s2_r[20] ), .CO(n551), .S0(n545) );
  HS65_GS_FA1X4 U617 ( .A0(n545), .B0(n544), .CI(n543), .CO(n550), .S0(n540)
         );
  HS65_GS_FA1X4 U618 ( .A0(n548), .B0(n547), .CI(n546), .CO(n553), .S0(n549)
         );
  HS65_GS_FA1X4 U619 ( .A0(n551), .B0(n550), .CI(n549), .CO(n1072), .S0(n1075)
         );
  HS65_GS_FA1X4 U620 ( .A0(n554), .B0(n553), .CI(n552), .CO(n1069), .S0(n1071)
         );
  HS65_GS_FA1X4 U621 ( .A0(n557), .B0(n556), .CI(n555), .CO(n1065), .S0(n1067)
         );
  HS65_GS_FA1X4 U622 ( .A0(\mul_b1/fa1_c1_r[22] ), .B0(\mul_b1/fa1_c2_r[22] ), 
        .CI(\mul_b1/fa1_s2_r[23] ), .CO(n563), .S0(n560) );
  HS65_GS_FA1X4 U623 ( .A0(n560), .B0(n559), .CI(n558), .CO(n562), .S0(n555)
         );
  HS65_GS_PAO2X4 U624 ( .A(\mul_b1/fa1_c0_r[22] ), .B(\mul_b1/fa1_s1_r[23] ), 
        .P(\mul_b1/fa1_s0_r[23] ), .Z(n565) );
  HS65_GSS_XOR3X2 U625 ( .A(\mul_b1/fa1_c0_r[23] ), .B(\mul_b1/fa1_s1_r[24] ), 
        .C(\mul_b1/fa1_s0_r[24] ), .Z(n564) );
  HS65_GS_FA1X4 U626 ( .A0(n563), .B0(n562), .CI(n561), .CO(n1060), .S0(n1063)
         );
  HS65_GS_FA1X4 U627 ( .A0(\mul_b1/fa1_c1_r[23] ), .B0(\mul_b1/fa1_c2_r[23] ), 
        .CI(\mul_b1/fa1_s2_r[24] ), .CO(n572), .S0(n566) );
  HS65_GS_FA1X4 U628 ( .A0(n566), .B0(n565), .CI(n564), .CO(n571), .S0(n561)
         );
  HS65_GS_FA1X4 U629 ( .A0(n569), .B0(n568), .CI(n567), .CO(n574), .S0(n570)
         );
  HS65_GS_FA1X4 U630 ( .A0(n572), .B0(n571), .CI(n570), .CO(n1056), .S0(n1059)
         );
  HS65_GS_FA1X4 U631 ( .A0(n575), .B0(n574), .CI(n573), .CO(n1053), .S0(n1055)
         );
  HS65_GS_FA1X4 U632 ( .A0(n578), .B0(n577), .CI(n576), .CO(n1030), .S0(n1051)
         );
  HS65_GS_FA1X4 U633 ( .A0(\mul_b1/fa1_c1_r[26] ), .B0(\mul_b1/fa1_c2_r[26] ), 
        .CI(\mul_b1/fa1_s2_r[27] ), .CO(n587), .S0(n581) );
  HS65_GS_FA1X4 U634 ( .A0(n581), .B0(n580), .CI(n579), .CO(n586), .S0(n576)
         );
  HS65_GS_FA1X4 U635 ( .A0(n584), .B0(n583), .CI(n582), .CO(n589), .S0(n585)
         );
  HS65_GS_FA1X4 U636 ( .A0(n587), .B0(n586), .CI(n585), .CO(n1035), .S0(n1028)
         );
  HS65_GS_FA1X4 U637 ( .A0(n590), .B0(n589), .CI(n588), .CO(n1033), .S0(n1034)
         );
  HS65_GS_FA1X4 U638 ( .A0(\mul_b1/fa1_c1_r[28] ), .B0(\mul_b1/fa1_c2_r[28] ), 
        .CI(\mul_b1/fa1_s2_r[29] ), .CO(n596), .S0(n593) );
  HS65_GS_FA1X4 U639 ( .A0(n593), .B0(n592), .CI(n591), .CO(n595), .S0(n588)
         );
  HS65_GS_PAO2X4 U640 ( .A(\mul_b1/fa1_c0_r[28] ), .B(\mul_b1/fa1_s1_r[29] ), 
        .P(\mul_b1/fa1_s0_r[29] ), .Z(n599) );
  HS65_GSS_XOR3X2 U641 ( .A(\mul_b1/fa1_c0_r[29] ), .B(\mul_b1/fa1_s1_r[30] ), 
        .C(\mul_b1/fa1_s0_r[30] ), .Z(n598) );
  HS65_GSS_XOR2X3 U642 ( .A(\mul_b1/fa1_s2_r[30] ), .B(\mul_b1/fa1_c1_r[29] ), 
        .Z(n597) );
  HS65_GS_FA1X4 U643 ( .A0(n596), .B0(n595), .CI(n594), .CO(n1041), .S0(n1031)
         );
  HS65_GS_AND2X4 U644 ( .A(\mul_b1/fa1_c1_r[29] ), .B(\mul_b1/fa1_s2_r[30] ), 
        .Z(n605) );
  HS65_GS_FA1X4 U645 ( .A0(n599), .B0(n598), .CI(n597), .CO(n604), .S0(n594)
         );
  HS65_GS_FA1X4 U646 ( .A0(n602), .B0(n601), .CI(n600), .CO(n414), .S0(n603)
         );
  HS65_GS_FA1X4 U647 ( .A0(n605), .B0(n604), .CI(n603), .CO(n1037), .S0(n1040)
         );
  HS65_GSS_XOR3X2 U648 ( .A(n606), .B(\mul_b1/fa1_s0_r[33] ), .C(
        \mul_b1/fa1_s2_r[33] ), .Z(n608) );
  HS65_GSS_XOR2X3 U649 ( .A(\mul_b1/fa1_c1_r[32] ), .B(\mul_b1/fa1_c0_r[32] ), 
        .Z(n607) );
  HS65_GSS_XOR3X2 U650 ( .A(n608), .B(\mul_b1/fa1_s1_r[33] ), .C(n607), .Z(
        n609) );
  HS65_GSS_XOR3X2 U651 ( .A(n611), .B(n610), .C(n609), .Z(n612) );
  HS65_GSS_XOR3X2 U652 ( .A(n614), .B(n613), .C(n612), .Z(
        \mul_b1/result_sat[15] ) );
  HS65_GS_IVX2 U653 ( .A(n1438), .Z(n1820) );
  HS65_GSS_XNOR2X3 U654 ( .A(n615), .B(n622), .Z(n629) );
  HS65_GS_FA1X4 U655 ( .A0(n618), .B0(n617), .CI(n616), .CO(n72), .S0(n628) );
  HS65_GS_FA1X4 U656 ( .A0(n621), .B0(n620), .CI(n619), .CO(n616), .S0(n627)
         );
  HS65_GS_AOI12X2 U657 ( .A(n624), .B(n623), .C(n622), .Z(n626) );
  HS65_GS_NAND3X2 U658 ( .A(n628), .B(n627), .C(n626), .Z(n625) );
  HS65_GS_OAI12X3 U659 ( .A(n629), .B(n625), .C(\mul_b0/result_sat[15] ), .Z(
        n1167) );
  HS65_GS_OAI21X2 U660 ( .A(n632), .B(n633), .C(n1167), .Z(n631) );
  HS65_GS_NOR3X1 U661 ( .A(n628), .B(n627), .C(n626), .Z(n630) );
  HS65_GS_AOI12X2 U662 ( .A(n630), .B(n629), .C(\mul_b0/result_sat[15] ), .Z(
        n1166) );
  HS65_GS_IVX2 U663 ( .A(n1166), .Z(n1806) );
  HS65_GS_CBI4I1X3 U664 ( .A(n633), .B(n632), .C(n631), .D(n1806), .Z(
        \mul_b0/result_sat[11] ) );
  HS65_GS_OAI21X2 U665 ( .A(n636), .B(n635), .C(n1167), .Z(n634) );
  HS65_GS_CBI4I1X3 U666 ( .A(n636), .B(n635), .C(n634), .D(n1806), .Z(
        \mul_b0/result_sat[5] ) );
  HS65_GS_NAND2X2 U667 ( .A(n639), .B(n638), .Z(n637) );
  HS65_GS_OAI21X2 U668 ( .A(n639), .B(n638), .C(n637), .Z(n643) );
  HS65_GS_IVX2 U669 ( .A(n640), .Z(n642) );
  HS65_GS_OAI21X2 U670 ( .A(n642), .B(n643), .C(n1167), .Z(n641) );
  HS65_GS_CBI4I1X3 U671 ( .A(n643), .B(n642), .C(n641), .D(n1806), .Z(
        \mul_b0/result_sat[4] ) );
  HS65_GS_OAI21X2 U672 ( .A(n646), .B(n645), .C(n644), .Z(n649) );
  HS65_GS_OAI21X2 U673 ( .A(n648), .B(n649), .C(n1167), .Z(n647) );
  HS65_GS_CBI4I1X3 U674 ( .A(n649), .B(n648), .C(n647), .D(n1806), .Z(
        \mul_b0/result_sat[2] ) );
  HS65_GSS_XOR2X3 U675 ( .A(x_z2[2]), .B(x_z2[4]), .Z(\mul_b1/fa1_s0[4] ) );
  HS65_GSS_XOR2X3 U676 ( .A(x_z2[1]), .B(x_z2[3]), .Z(\mul_b1/fa1_s0[3] ) );
  HS65_GS_IVX2 U677 ( .A(x_z2[14]), .Z(n1745) );
  HS65_GS_IVX2 U678 ( .A(x_z2[11]), .Z(n1432) );
  HS65_GS_IVX2 U679 ( .A(x_z2[10]), .Z(n1429) );
  HS65_GS_IVX2 U680 ( .A(x_z2[9]), .Z(n1428) );
  HS65_GS_IVX2 U681 ( .A(x_z2[7]), .Z(n1423) );
  HS65_GS_IVX2 U682 ( .A(x_z2[6]), .Z(n1421) );
  HS65_GS_IVX2 U683 ( .A(x_z2[5]), .Z(n1419) );
  HS65_GS_IVX2 U684 ( .A(x_z2[4]), .Z(n1418) );
  HS65_GS_IVX2 U685 ( .A(x_z2[3]), .Z(n1416) );
  HS65_GS_IVX2 U686 ( .A(x_z2[2]), .Z(n1414) );
  HS65_GS_IVX2 U687 ( .A(x_z2[1]), .Z(n1752) );
  HS65_GS_IVX2 U688 ( .A(y_z2[14]), .Z(n1676) );
  HS65_GS_IVX2 U689 ( .A(y_z2[13]), .Z(n1678) );
  HS65_GS_IVX2 U690 ( .A(y_z2[12]), .Z(n1680) );
  HS65_GS_IVX2 U691 ( .A(y_z2[11]), .Z(n1682) );
  HS65_GS_IVX2 U692 ( .A(y_z2[10]), .Z(n1684) );
  HS65_GS_IVX2 U693 ( .A(y_z2[9]), .Z(n1686) );
  HS65_GS_IVX2 U694 ( .A(y_z2[8]), .Z(n1688) );
  HS65_GS_IVX2 U695 ( .A(y_z2[7]), .Z(n1690) );
  HS65_GS_IVX2 U696 ( .A(y_z2[6]), .Z(n1692) );
  HS65_GS_IVX2 U697 ( .A(y_z2[5]), .Z(n1694) );
  HS65_GS_IVX2 U698 ( .A(y_z2[4]), .Z(n1696) );
  HS65_GS_IVX2 U699 ( .A(y_z2[3]), .Z(n1698) );
  HS65_GS_IVX2 U700 ( .A(y_z2[2]), .Z(n1700) );
  HS65_GS_IVX2 U701 ( .A(y_z2[1]), .Z(n1702) );
  HS65_GS_IVX2 U702 ( .A(y_z2[0]), .Z(n1701) );
  HS65_GS_NOR2X2 U703 ( .A(y_z2[15]), .B(n1674), .Z(n1814) );
  HS65_GSS_XNOR2X3 U704 ( .A(n650), .B(n657), .Z(n664) );
  HS65_GS_FA1X4 U705 ( .A0(n653), .B0(n652), .CI(n651), .CO(n170), .S0(n663)
         );
  HS65_GS_FA1X4 U706 ( .A0(n656), .B0(n655), .CI(n654), .CO(n651), .S0(n662)
         );
  HS65_GS_AOI12X2 U707 ( .A(n659), .B(n658), .C(n657), .Z(n661) );
  HS65_GS_NAND3X2 U708 ( .A(n663), .B(n662), .C(n661), .Z(n660) );
  HS65_GS_OAI12X3 U709 ( .A(n664), .B(n660), .C(\mul_a2/result_sat[15] ), .Z(
        n1341) );
  HS65_GS_OAI21X2 U710 ( .A(n667), .B(n668), .C(n1341), .Z(n666) );
  HS65_GS_NOR3X1 U711 ( .A(n663), .B(n662), .C(n661), .Z(n665) );
  HS65_GS_AOI12X2 U712 ( .A(n665), .B(n664), .C(\mul_a2/result_sat[15] ), .Z(
        n1340) );
  HS65_GS_IVX2 U713 ( .A(n1340), .Z(n1763) );
  HS65_GS_CBI4I1X3 U714 ( .A(n668), .B(n667), .C(n666), .D(n1763), .Z(
        \mul_a2/result_sat[14] ) );
  HS65_GSS_XOR2X3 U715 ( .A(n670), .B(n669), .Z(n673) );
  HS65_GS_OAI21X2 U716 ( .A(n672), .B(n673), .C(n1341), .Z(n671) );
  HS65_GS_CBI4I1X3 U717 ( .A(n673), .B(n672), .C(n671), .D(n1763), .Z(
        \mul_a2/result_sat[13] ) );
  HS65_GS_OAI21X2 U718 ( .A(n676), .B(n675), .C(n1341), .Z(n674) );
  HS65_GS_CBI4I1X3 U719 ( .A(n676), .B(n675), .C(n674), .D(n1763), .Z(
        \mul_a2/result_sat[5] ) );
  HS65_GS_NAND2X2 U720 ( .A(n679), .B(n678), .Z(n677) );
  HS65_GS_OAI21X2 U721 ( .A(n679), .B(n678), .C(n677), .Z(n683) );
  HS65_GS_IVX2 U722 ( .A(n680), .Z(n682) );
  HS65_GS_OAI21X2 U723 ( .A(n682), .B(n683), .C(n1341), .Z(n681) );
  HS65_GS_CBI4I1X3 U724 ( .A(n683), .B(n682), .C(n681), .D(n1763), .Z(
        \mul_a2/result_sat[4] ) );
  HS65_GS_OAI21X2 U725 ( .A(n686), .B(n685), .C(n684), .Z(n689) );
  HS65_GS_OAI21X2 U726 ( .A(n688), .B(n689), .C(n1341), .Z(n687) );
  HS65_GS_CBI4I1X3 U727 ( .A(n689), .B(n688), .C(n687), .D(n1763), .Z(
        \mul_a2/result_sat[2] ) );
  HS65_GS_IVX2 U728 ( .A(y_z1[14]), .Z(n1724) );
  HS65_GS_IVX2 U729 ( .A(y_z1[13]), .Z(n1726) );
  HS65_GS_IVX2 U730 ( .A(y_z1[12]), .Z(n1728) );
  HS65_GS_IVX2 U731 ( .A(y_z1[11]), .Z(n1730) );
  HS65_GS_IVX2 U732 ( .A(y_z1[10]), .Z(n1732) );
  HS65_GS_IVX2 U733 ( .A(y_z1[9]), .Z(n1734) );
  HS65_GS_IVX2 U734 ( .A(y_z1[8]), .Z(n1736) );
  HS65_GS_IVX2 U735 ( .A(y_z1[7]), .Z(n1738) );
  HS65_GS_IVX2 U736 ( .A(y_z1[6]), .Z(n1740) );
  HS65_GS_IVX2 U737 ( .A(y_z1[5]), .Z(n1716) );
  HS65_GS_IVX2 U738 ( .A(y_z1[4]), .Z(n1718) );
  HS65_GS_IVX2 U739 ( .A(y_z1[3]), .Z(n1720) );
  HS65_GS_IVX2 U740 ( .A(y_z1[2]), .Z(n1754) );
  HS65_GS_IVX2 U741 ( .A(y_z1[1]), .Z(n1755) );
  HS65_GS_IVX2 U742 ( .A(\mul_a1/fa1_s1[7] ), .Z(n1753) );
  HS65_GS_HA1X4 U743 ( .A0(n1755), .B0(n1753), .CO(n690) );
  HS65_GS_HA1X4 U744 ( .A0(n1754), .B0(n690), .CO(n691) );
  HS65_GS_HA1X4 U745 ( .A0(n1720), .B0(n691), .CO(n692) );
  HS65_GS_HA1X4 U746 ( .A0(n1718), .B0(n692), .CO(n693) );
  HS65_GS_HA1X4 U747 ( .A0(n1716), .B0(n693), .CO(n1739) );
  HS65_GS_NOR2X5 U748 ( .A(n1819), .B(n1722), .Z(n1811) );
  HS65_GS_IVX2 U749 ( .A(n1705), .Z(n1819) );
  HS65_GS_BFX4 U750 ( .A(valid_in), .Z(n1440) );
  HS65_GS_MUX21I1X3 U751 ( .D0(n1754), .D1(data_out[2]), .S0(n1440), .Z(n1910)
         );
  HS65_GS_MUX21I1X3 U752 ( .D0(n1720), .D1(data_out[3]), .S0(n1440), .Z(n1907)
         );
  HS65_GS_MUX21I1X3 U753 ( .D0(n1740), .D1(data_out[6]), .S0(n1440), .Z(n1898)
         );
  HS65_GS_MUX21I1X3 U754 ( .D0(n1738), .D1(data_out[7]), .S0(n1440), .Z(n1895)
         );
  HS65_GS_AND2X4 U755 ( .A(p_b1[1]), .B(p_b0[1]), .Z(n705) );
  HS65_GSS_XOR2X3 U756 ( .A(p_b1[1]), .B(p_b0[1]), .Z(n708) );
  HS65_GS_FA1X4 U757 ( .A0(p_b0[2]), .B0(p_b1[2]), .CI(p_b2[2]), .CO(n701), 
        .S0(n703) );
  HS65_GS_FA1X4 U758 ( .A0(p_b0[3]), .B0(p_b1[3]), .CI(p_b2[3]), .CO(n722), 
        .S0(n699) );
  HS65_GS_FA1X4 U759 ( .A0(p_b0[4]), .B0(p_b1[4]), .CI(p_b2[4]), .CO(n697), 
        .S0(n720) );
  HS65_GS_FA1X4 U760 ( .A0(p_b0[5]), .B0(p_b1[5]), .CI(p_b2[5]), .CO(n731), 
        .S0(n695) );
  HS65_GS_IVX2 U761 ( .A(n694), .Z(n728) );
  HS65_GS_FA1X4 U762 ( .A0(n697), .B0(n696), .CI(n695), .CO(n730), .S0(n698)
         );
  HS65_GS_IVX2 U763 ( .A(n698), .Z(n727) );
  HS65_GS_FA1X4 U764 ( .A0(n701), .B0(n700), .CI(n699), .CO(n721), .S0(n702)
         );
  HS65_GS_IVX2 U765 ( .A(n702), .Z(n716) );
  HS65_GS_FA1X4 U766 ( .A0(n705), .B0(n704), .CI(n703), .CO(n700), .S0(n706)
         );
  HS65_GS_IVX2 U767 ( .A(n706), .Z(n711) );
  HS65_GS_FA1X4 U768 ( .A0(p_b2[1]), .B0(n708), .CI(n707), .CO(n704), .S0(n709) );
  HS65_GS_IVX2 U769 ( .A(n709), .Z(n713) );
  HS65_GS_FA1X4 U770 ( .A0(p_b2[0]), .B0(p_b0[0]), .CI(p_b1[0]), .CO(n707), 
        .S0(n710) );
  HS65_GS_IVX2 U771 ( .A(n710), .Z(n1444) );
  HS65_GS_NAND2X2 U772 ( .A(n1350), .B(p_a1[1]), .Z(n1349) );
  HS65_GS_NAND3AX3 U773 ( .A(n1349), .B(p_a2[1]), .C(n713), .Z(n715) );
  HS65_GS_FA1X4 U774 ( .A0(p_a2[2]), .B0(p_a1[2]), .CI(n711), .CO(n718), .S0(
        n1354) );
  HS65_GS_FA1X4 U775 ( .A0(p_a2[1]), .B0(n713), .CI(n712), .CO(n714), .S0(
        n1350) );
  HS65_GS_CB4I1X4 U776 ( .A(p_a1[1]), .B(n1350), .C(n714), .D(n715), .Z(n1353)
         );
  HS65_GS_NAND2X2 U777 ( .A(n1354), .B(n1353), .Z(n1352) );
  HS65_GS_NAND2X2 U778 ( .A(n715), .B(n1352), .Z(n717) );
  HS65_GS_NOR2X2 U779 ( .A(n718), .B(n717), .Z(n719) );
  HS65_GS_FA1X4 U780 ( .A0(p_a2[3]), .B0(p_a1[3]), .CI(n716), .CO(n1361), .S0(
        n1358) );
  HS65_GSS_XNOR2X3 U781 ( .A(n718), .B(n717), .Z(n1357) );
  HS65_GS_NOR2X2 U782 ( .A(n1358), .B(n1357), .Z(n1356) );
  HS65_GS_NOR2X2 U783 ( .A(n719), .B(n1356), .Z(n1360) );
  HS65_GS_FA1X4 U784 ( .A0(n722), .B0(n721), .CI(n720), .CO(n696), .S0(n723)
         );
  HS65_GS_IVX2 U785 ( .A(n723), .Z(n724) );
  HS65_GS_PAO2X4 U786 ( .A(n1361), .B(n1360), .P(n1363), .Z(n725) );
  HS65_GS_FA1X4 U787 ( .A0(p_a2[4]), .B0(p_a1[4]), .CI(n724), .CO(n726), .S0(
        n1363) );
  HS65_GSS_XOR2X3 U788 ( .A(n725), .B(n726), .Z(n1369) );
  HS65_GS_AO22X4 U789 ( .A(n1368), .B(n1369), .C(n726), .D(n725), .Z(n1374) );
  HS65_GS_FA1X4 U790 ( .A0(p_a2[5]), .B0(p_a1[5]), .CI(n727), .CO(n1373), .S0(
        n1368) );
  HS65_GS_FA1X4 U791 ( .A0(p_a2[6]), .B0(p_a1[6]), .CI(n728), .CO(n767), .S0(
        n1372) );
  HS65_GS_FA1X4 U792 ( .A0(p_b0[6]), .B0(p_b1[6]), .CI(p_b2[6]), .CO(n735), 
        .S0(n729) );
  HS65_GS_FA1X4 U793 ( .A0(n731), .B0(n730), .CI(n729), .CO(n734), .S0(n694)
         );
  HS65_GS_IVX2 U794 ( .A(n732), .Z(n768) );
  HS65_GS_FA1X4 U795 ( .A0(p_b0[7]), .B0(p_b1[7]), .CI(p_b2[7]), .CO(n763), 
        .S0(n733) );
  HS65_GS_FA1X4 U796 ( .A0(n735), .B0(n734), .CI(n733), .CO(n762), .S0(n732)
         );
  HS65_GS_FA1X4 U797 ( .A0(p_b0[8]), .B0(p_b1[8]), .CI(p_b2[8]), .CO(n759), 
        .S0(n761) );
  HS65_GS_FA1X4 U798 ( .A0(p_b0[9]), .B0(p_b1[9]), .CI(p_b2[9]), .CO(n755), 
        .S0(n757) );
  HS65_GS_FA1X4 U799 ( .A0(p_b0[10]), .B0(p_b1[10]), .CI(p_b2[10]), .CO(n751), 
        .S0(n753) );
  HS65_GS_FA1X4 U800 ( .A0(p_b0[11]), .B0(p_b1[11]), .CI(p_b2[11]), .CO(n743), 
        .S0(n749) );
  HS65_GS_FA1X4 U801 ( .A0(p_b0[12]), .B0(p_b1[12]), .CI(p_b2[12]), .CO(n747), 
        .S0(n741) );
  HS65_GS_FA1X4 U802 ( .A0(p_b0[13]), .B0(p_b1[13]), .CI(p_b2[13]), .CO(n739), 
        .S0(n745) );
  HS65_GS_FA1X4 U803 ( .A0(p_b0[14]), .B0(p_b1[14]), .CI(p_b2[14]), .CO(n791), 
        .S0(n737) );
  HS65_GS_IVX2 U804 ( .A(p_b0[15]), .Z(n792) );
  HS65_GS_NAND2X2 U805 ( .A(p_b2[15]), .B(p_b1[15]), .Z(n793) );
  HS65_GS_OAI21X2 U806 ( .A(p_b2[15]), .B(p_b1[15]), .C(n793), .Z(n736) );
  HS65_GS_MUXI21X2 U807 ( .D0(p_b0[15]), .D1(n792), .S0(n736), .Z(n789) );
  HS65_GS_FA1X4 U808 ( .A0(n739), .B0(n738), .CI(n737), .CO(n790), .S0(n740)
         );
  HS65_GS_IVX2 U809 ( .A(n740), .Z(n786) );
  HS65_GS_FA1X4 U810 ( .A0(n743), .B0(n742), .CI(n741), .CO(n746), .S0(n744)
         );
  HS65_GS_IVX2 U811 ( .A(n744), .Z(n779) );
  HS65_GS_FA1X4 U812 ( .A0(n747), .B0(n746), .CI(n745), .CO(n738), .S0(n748)
         );
  HS65_GS_IVX2 U813 ( .A(n748), .Z(n783) );
  HS65_GS_FA1X4 U814 ( .A0(n751), .B0(n750), .CI(n749), .CO(n742), .S0(n752)
         );
  HS65_GS_IVX2 U815 ( .A(n752), .Z(n775) );
  HS65_GS_FA1X4 U816 ( .A0(n755), .B0(n754), .CI(n753), .CO(n750), .S0(n756)
         );
  HS65_GS_IVX2 U817 ( .A(n756), .Z(n771) );
  HS65_GS_FA1X4 U818 ( .A0(n759), .B0(n758), .CI(n757), .CO(n754), .S0(n760)
         );
  HS65_GS_IVX2 U819 ( .A(n760), .Z(n770) );
  HS65_GS_FA1X4 U820 ( .A0(n763), .B0(n762), .CI(n761), .CO(n758), .S0(n764)
         );
  HS65_GS_IVX2 U821 ( .A(n764), .Z(n769) );
  HS65_GS_FA1X4 U822 ( .A0(n767), .B0(n766), .CI(n765), .CO(n813), .S0(n810)
         );
  HS65_GS_FA1X4 U823 ( .A0(p_a2[7]), .B0(p_a1[7]), .CI(n768), .CO(n812), .S0(
        n765) );
  HS65_GS_FA1X4 U824 ( .A0(p_a2[8]), .B0(p_a1[8]), .CI(n769), .CO(n1378), .S0(
        n811) );
  HS65_GS_FA1X4 U825 ( .A0(p_a2[9]), .B0(p_a1[9]), .CI(n770), .CO(n772), .S0(
        n1380) );
  HS65_GS_PAO2X4 U826 ( .A(n1378), .B(n1377), .P(n1380), .Z(n773) );
  HS65_GS_NAND2X2 U827 ( .A(n772), .B(n773), .Z(n774) );
  HS65_GS_FA1X4 U828 ( .A0(p_a2[10]), .B0(p_a1[10]), .CI(n771), .CO(n776), 
        .S0(n1386) );
  HS65_GSS_XOR2X3 U829 ( .A(n773), .B(n772), .Z(n1385) );
  HS65_GS_NAND2X2 U830 ( .A(n1386), .B(n1385), .Z(n1384) );
  HS65_GS_NAND2X2 U831 ( .A(n774), .B(n1384), .Z(n777) );
  HS65_GS_NAND2X2 U832 ( .A(n776), .B(n777), .Z(n778) );
  HS65_GS_FA1X4 U833 ( .A0(p_a2[11]), .B0(p_a1[11]), .CI(n775), .CO(n780), 
        .S0(n1390) );
  HS65_GSS_XOR2X3 U834 ( .A(n777), .B(n776), .Z(n1389) );
  HS65_GS_NAND2X2 U835 ( .A(n1390), .B(n1389), .Z(n1388) );
  HS65_GS_NAND2X2 U836 ( .A(n778), .B(n1388), .Z(n781) );
  HS65_GS_NAND2X2 U837 ( .A(n780), .B(n781), .Z(n782) );
  HS65_GS_FA1X4 U838 ( .A0(p_a2[12]), .B0(p_a1[12]), .CI(n779), .CO(n1396), 
        .S0(n1394) );
  HS65_GSS_XOR2X3 U839 ( .A(n781), .B(n780), .Z(n1393) );
  HS65_GS_NAND2X2 U840 ( .A(n1394), .B(n1393), .Z(n1392) );
  HS65_GS_NAND2X2 U841 ( .A(n782), .B(n1392), .Z(n1397) );
  HS65_GS_PAO2X4 U842 ( .A(n1396), .B(n1399), .P(n1397), .Z(n784) );
  HS65_GS_FA1X4 U843 ( .A0(p_a1[13]), .B0(p_a2[13]), .CI(n783), .CO(n785), 
        .S0(n1399) );
  HS65_GSS_XOR2X3 U844 ( .A(n784), .B(n785), .Z(n1407) );
  HS65_GS_AO22X4 U845 ( .A(n1406), .B(n1407), .C(n785), .D(n784), .Z(n798) );
  HS65_GS_FA1X4 U846 ( .A0(p_a1[14]), .B0(p_a2[14]), .CI(n786), .CO(n797), 
        .S0(n1406) );
  HS65_GS_FA1X4 U847 ( .A0(p_a1[15]), .B0(p_a2[15]), .CI(n787), .CO(n803), 
        .S0(n788) );
  HS65_GS_IVX2 U848 ( .A(n788), .Z(n796) );
  HS65_GS_FA1X4 U849 ( .A0(n791), .B0(n790), .CI(n789), .CO(n795), .S0(n787)
         );
  HS65_GS_OAI32X2 U850 ( .A(p_b0[15]), .B(p_b2[15]), .C(p_b1[15]), .D(n793), 
        .E(n792), .Z(n794) );
  HS65_GSS_XNOR2X3 U851 ( .A(n795), .B(n794), .Z(n800) );
  HS65_GSS_XNOR2X3 U852 ( .A(n801), .B(n800), .Z(n802) );
  HS65_GS_AND2X4 U853 ( .A(n803), .B(n802), .Z(n805) );
  HS65_GS_FA1X4 U854 ( .A0(n798), .B0(n797), .CI(n796), .CO(n801), .S0(n799)
         );
  HS65_GS_IVX2 U855 ( .A(n799), .Z(n808) );
  HS65_GS_NAND2X2 U856 ( .A(n801), .B(n800), .Z(n804) );
  HS65_GS_IVX2 U857 ( .A(valid_T3), .Z(n1810) );
  HS65_GS_NOR2X2 U858 ( .A(n803), .B(n802), .Z(n806) );
  HS65_GS_NOR3AX2 U859 ( .A(n804), .B(n1810), .C(n806), .Z(n1808) );
  HS65_GS_OAI12X3 U860 ( .A(n805), .B(n808), .C(n1808), .Z(n1403) );
  HS65_GS_OA12X4 U861 ( .A(n806), .B(n805), .C(valid_T3), .Z(n807) );
  HS65_GS_AOI12X2 U862 ( .A(n808), .B(n807), .C(n1808), .Z(n1448) );
  HS65_GS_NAND2X2 U863 ( .A(data_out[7]), .B(n1810), .Z(n809) );
  HS65_GS_CBI4I1X3 U864 ( .A(n810), .B(n1403), .C(n1448), .D(n809), .Z(n1894)
         );
  HS65_GS_MUX21I1X3 U865 ( .D0(n1736), .D1(data_out[8]), .S0(n1440), .Z(n1892)
         );
  HS65_GS_FA1X4 U866 ( .A0(n813), .B0(n812), .CI(n811), .CO(n1377), .S0(n815)
         );
  HS65_GS_NAND2X2 U867 ( .A(data_out[8]), .B(n1810), .Z(n814) );
  HS65_GS_CBI4I1X3 U868 ( .A(n815), .B(n1403), .C(n1448), .D(n814), .Z(n1891)
         );
  HS65_GS_MUX21I1X3 U869 ( .D0(n1732), .D1(data_out[10]), .S0(n1440), .Z(n1886) );
  HS65_GS_MUX21I1X3 U870 ( .D0(n1730), .D1(data_out[11]), .S0(n1440), .Z(n1883) );
  HS65_GS_MUX21I1X3 U871 ( .D0(n1728), .D1(data_out[12]), .S0(n1440), .Z(n1880) );
  HS65_GSS_XNOR2X3 U872 ( .A(n817), .B(n816), .Z(n839) );
  HS65_GS_IVX2 U873 ( .A(n818), .Z(n838) );
  HS65_GS_FA1X4 U874 ( .A0(n821), .B0(n820), .CI(n819), .CO(n823), .S0(n836)
         );
  HS65_GS_FA1X4 U875 ( .A0(n824), .B0(n823), .CI(n822), .CO(n829), .S0(n834)
         );
  HS65_GS_FA1X4 U876 ( .A0(n827), .B0(n826), .CI(n825), .CO(n820), .S0(n833)
         );
  HS65_GS_FA1X4 U877 ( .A0(n830), .B0(n829), .CI(n828), .CO(n402), .S0(n832)
         );
  HS65_GS_OR3X4 U878 ( .A(n834), .B(n833), .C(n832), .Z(n831) );
  HS65_GS_OAI21X2 U879 ( .A(n836), .B(n831), .C(\mul_b2/result_sat[15] ), .Z(
        n1571) );
  HS65_GS_OAI21X2 U880 ( .A(n838), .B(n839), .C(n1571), .Z(n837) );
  HS65_GS_AND3X4 U881 ( .A(n834), .B(n833), .C(n832), .Z(n835) );
  HS65_GS_AOI12X2 U882 ( .A(n836), .B(n835), .C(\mul_b2/result_sat[15] ), .Z(
        n1570) );
  HS65_GS_IVX2 U883 ( .A(n1570), .Z(n1791) );
  HS65_GS_CBI4I1X3 U884 ( .A(n839), .B(n838), .C(n837), .D(n1791), .Z(
        \mul_b2/result_sat[12] ) );
  HS65_GSS_XNOR2X3 U885 ( .A(n841), .B(n840), .Z(n844) );
  HS65_GS_OAI21X2 U886 ( .A(n843), .B(n844), .C(n1571), .Z(n842) );
  HS65_GS_CBI4I1X3 U887 ( .A(n844), .B(n843), .C(n842), .D(n1791), .Z(
        \mul_b2/result_sat[7] ) );
  HS65_GS_OAI21X2 U888 ( .A(n846), .B(n847), .C(n1571), .Z(n845) );
  HS65_GS_CBI4I1X3 U889 ( .A(n847), .B(n846), .C(n845), .D(n1791), .Z(
        \mul_b2/result_sat[2] ) );
  HS65_GS_IVX2 U890 ( .A(x_z2[13]), .Z(n1747) );
  HS65_GS_IVX2 U891 ( .A(x_z2[12]), .Z(n1749) );
  HS65_GS_IVX2 U892 ( .A(x_z2[8]), .Z(n1425) );
  HS65_GS_NOR2X3 U893 ( .A(\DP_OP_331J1_157_5454/n87 ), .B(n1743), .Z(n1813)
         );
  HS65_GS_NOR2X2 U894 ( .A(n1755), .B(n1754), .Z(\mul_a1/fa1_c1[9] ) );
  HS65_GS_NOR2X2 U895 ( .A(n1753), .B(n1755), .Z(\mul_a1/fa1_c1[8] ) );
  HS65_GS_NOR2X2 U896 ( .A(y_z1[15]), .B(n1703), .Z(n1815) );
  HS65_GS_AND2X4 U897 ( .A(\mul_a1/fa1_s2_r[31] ), .B(\mul_a1/fa1_c1_r[30] ), 
        .Z(n1003) );
  HS65_GS_AND2X4 U898 ( .A(\mul_a1/fa1_s1_r[31] ), .B(\mul_a1/fa1_s0_r[31] ), 
        .Z(n1006) );
  HS65_GSS_XOR2X3 U899 ( .A(\mul_a1/fa1_s2_r[32] ), .B(\mul_a1/fa1_c1_r[31] ), 
        .Z(n1005) );
  HS65_GS_NAND2X2 U900 ( .A(\mul_a1/fa1_s1_r[32] ), .B(\mul_a1/fa1_s0_r[32] ), 
        .Z(n1007) );
  HS65_GS_OA12X4 U901 ( .A(\mul_a1/fa1_s1_r[32] ), .B(\mul_a1/fa1_s0_r[32] ), 
        .C(n1007), .Z(n1004) );
  HS65_GSS_XOR2X3 U902 ( .A(\mul_a1/fa1_s2_r[31] ), .B(\mul_a1/fa1_c1_r[30] ), 
        .Z(n994) );
  HS65_GSS_XOR2X3 U903 ( .A(\mul_a1/fa1_s1_r[31] ), .B(\mul_a1/fa1_s0_r[31] ), 
        .Z(n993) );
  HS65_GS_AND2X4 U904 ( .A(\mul_a1/fa1_s0_r[30] ), .B(\mul_a1/fa1_s1_r[30] ), 
        .Z(n992) );
  HS65_GS_AND2X4 U905 ( .A(\mul_a1/fa1_s2_r[29] ), .B(\mul_a1/fa1_c1_r[28] ), 
        .Z(n991) );
  HS65_GSS_XOR2X3 U906 ( .A(\mul_a1/fa1_s2_r[29] ), .B(\mul_a1/fa1_c1_r[28] ), 
        .Z(n850) );
  HS65_GSS_XOR2X3 U907 ( .A(\mul_a1/fa1_s1_r[29] ), .B(\mul_a1/fa1_s0_r[29] ), 
        .Z(n849) );
  HS65_GS_AND2X4 U908 ( .A(\mul_a1/fa1_s0_r[28] ), .B(\mul_a1/fa1_s1_r[28] ), 
        .Z(n848) );
  HS65_GS_AND2X4 U909 ( .A(\mul_a1/fa1_s1_r[29] ), .B(\mul_a1/fa1_s0_r[29] ), 
        .Z(n997) );
  HS65_GSS_XOR2X3 U910 ( .A(\mul_a1/fa1_s2_r[30] ), .B(\mul_a1/fa1_c1_r[29] ), 
        .Z(n996) );
  HS65_GSS_XOR2X3 U911 ( .A(\mul_a1/fa1_s0_r[30] ), .B(\mul_a1/fa1_s1_r[30] ), 
        .Z(n995) );
  HS65_GS_AND2X4 U912 ( .A(\mul_a1/fa1_s2_r[28] ), .B(\mul_a1/fa1_c1_r[27] ), 
        .Z(n988) );
  HS65_GSS_XOR2X3 U913 ( .A(\mul_a1/fa1_s2_r[28] ), .B(\mul_a1/fa1_c1_r[27] ), 
        .Z(n982) );
  HS65_GSS_XOR2X3 U914 ( .A(\mul_a1/fa1_s0_r[28] ), .B(\mul_a1/fa1_s1_r[28] ), 
        .Z(n981) );
  HS65_GS_AND2X4 U915 ( .A(\mul_a1/fa1_s1_r[27] ), .B(\mul_a1/fa1_s0_r[27] ), 
        .Z(n980) );
  HS65_GS_FA1X4 U916 ( .A0(n850), .B0(n849), .CI(n848), .CO(n990), .S0(n986)
         );
  HS65_GS_AND2X4 U917 ( .A(\mul_a1/fa1_s2_r[26] ), .B(\mul_a1/fa1_c1_r[25] ), 
        .Z(n976) );
  HS65_GSS_XOR2X3 U918 ( .A(\mul_a1/fa1_s2_r[26] ), .B(\mul_a1/fa1_c1_r[25] ), 
        .Z(n853) );
  HS65_GSS_XOR2X3 U919 ( .A(\mul_a1/fa1_s1_r[26] ), .B(\mul_a1/fa1_s0_r[26] ), 
        .Z(n852) );
  HS65_GS_AND2X4 U920 ( .A(\mul_a1/fa1_s0_r[25] ), .B(\mul_a1/fa1_s1_r[25] ), 
        .Z(n851) );
  HS65_GS_AND2X4 U921 ( .A(\mul_a1/fa1_s1_r[26] ), .B(\mul_a1/fa1_s0_r[26] ), 
        .Z(n979) );
  HS65_GSS_XOR2X3 U922 ( .A(\mul_a1/fa1_s2_r[27] ), .B(\mul_a1/fa1_c1_r[26] ), 
        .Z(n978) );
  HS65_GSS_XOR2X3 U923 ( .A(\mul_a1/fa1_s1_r[27] ), .B(\mul_a1/fa1_s0_r[27] ), 
        .Z(n977) );
  HS65_GS_AND2X4 U924 ( .A(\mul_a1/fa1_s2_r[25] ), .B(\mul_a1/fa1_c1_r[24] ), 
        .Z(n973) );
  HS65_GSS_XOR2X3 U925 ( .A(\mul_a1/fa1_s2_r[25] ), .B(\mul_a1/fa1_c1_r[24] ), 
        .Z(n856) );
  HS65_GSS_XOR2X3 U926 ( .A(\mul_a1/fa1_s0_r[25] ), .B(\mul_a1/fa1_s1_r[25] ), 
        .Z(n855) );
  HS65_GS_AND2X4 U927 ( .A(\mul_a1/fa1_s0_r[24] ), .B(\mul_a1/fa1_s1_r[24] ), 
        .Z(n854) );
  HS65_GS_FA1X4 U928 ( .A0(n853), .B0(n852), .CI(n851), .CO(n975), .S0(n971)
         );
  HS65_GS_AND2X4 U929 ( .A(\mul_a1/fa1_s2_r[24] ), .B(\mul_a1/fa1_c1_r[23] ), 
        .Z(n970) );
  HS65_GSS_XOR2X3 U930 ( .A(\mul_a1/fa1_s2_r[24] ), .B(\mul_a1/fa1_c1_r[23] ), 
        .Z(n964) );
  HS65_GSS_XOR2X3 U931 ( .A(\mul_a1/fa1_s0_r[24] ), .B(\mul_a1/fa1_s1_r[24] ), 
        .Z(n963) );
  HS65_GS_AND2X4 U932 ( .A(\mul_a1/fa1_s1_r[23] ), .B(\mul_a1/fa1_s0_r[23] ), 
        .Z(n962) );
  HS65_GS_FA1X4 U933 ( .A0(n856), .B0(n855), .CI(n854), .CO(n972), .S0(n968)
         );
  HS65_GS_AND2X4 U934 ( .A(\mul_a1/fa1_s2_r[22] ), .B(\mul_a1/fa1_c1_r[21] ), 
        .Z(n958) );
  HS65_GSS_XOR2X3 U935 ( .A(\mul_a1/fa1_s2_r[22] ), .B(\mul_a1/fa1_c1_r[21] ), 
        .Z(n952) );
  HS65_GSS_XOR2X3 U936 ( .A(\mul_a1/fa1_s1_r[22] ), .B(\mul_a1/fa1_s0_r[22] ), 
        .Z(n951) );
  HS65_GS_AND2X4 U937 ( .A(\mul_a1/fa1_s1_r[21] ), .B(\mul_a1/fa1_s0_r[21] ), 
        .Z(n950) );
  HS65_GS_AND2X4 U938 ( .A(\mul_a1/fa1_s1_r[22] ), .B(\mul_a1/fa1_s0_r[22] ), 
        .Z(n961) );
  HS65_GSS_XOR2X3 U939 ( .A(\mul_a1/fa1_s2_r[23] ), .B(\mul_a1/fa1_c1_r[22] ), 
        .Z(n960) );
  HS65_GSS_XOR2X3 U940 ( .A(\mul_a1/fa1_s1_r[23] ), .B(\mul_a1/fa1_s0_r[23] ), 
        .Z(n959) );
  HS65_GS_AND2X4 U941 ( .A(\mul_a1/fa1_s2_r[20] ), .B(\mul_a1/fa1_c1_r[19] ), 
        .Z(n946) );
  HS65_GSS_XOR2X3 U942 ( .A(\mul_a1/fa1_s2_r[20] ), .B(\mul_a1/fa1_c1_r[19] ), 
        .Z(n859) );
  HS65_GSS_XOR2X3 U943 ( .A(\mul_a1/fa1_s1_r[20] ), .B(\mul_a1/fa1_s0_r[20] ), 
        .Z(n858) );
  HS65_GS_AND2X4 U944 ( .A(\mul_a1/fa1_s0_r[19] ), .B(\mul_a1/fa1_s1_r[19] ), 
        .Z(n857) );
  HS65_GS_AND2X4 U945 ( .A(\mul_a1/fa1_s1_r[20] ), .B(\mul_a1/fa1_s0_r[20] ), 
        .Z(n949) );
  HS65_GSS_XOR2X3 U946 ( .A(\mul_a1/fa1_s2_r[21] ), .B(\mul_a1/fa1_c1_r[20] ), 
        .Z(n948) );
  HS65_GSS_XOR2X3 U947 ( .A(\mul_a1/fa1_s1_r[21] ), .B(\mul_a1/fa1_s0_r[21] ), 
        .Z(n947) );
  HS65_GS_AND2X4 U948 ( .A(\mul_a1/fa1_c1_r[18] ), .B(\mul_a1/fa1_s2_r[19] ), 
        .Z(n862) );
  HS65_GSS_XOR2X3 U949 ( .A(\mul_a1/fa1_s0_r[19] ), .B(\mul_a1/fa1_s1_r[19] ), 
        .Z(n940) );
  HS65_GSS_XOR2X3 U950 ( .A(\mul_a1/fa1_c1_r[18] ), .B(\mul_a1/fa1_s2_r[19] ), 
        .Z(n939) );
  HS65_GS_AND2X4 U951 ( .A(\mul_a1/fa1_s1_r[18] ), .B(\mul_a1/fa1_s0_r[18] ), 
        .Z(n938) );
  HS65_GS_FA1X4 U952 ( .A0(n859), .B0(n858), .CI(n857), .CO(n945), .S0(n860)
         );
  HS65_GS_FA1X4 U953 ( .A0(n862), .B0(n861), .CI(n860), .CO(n1645), .S0(n1652)
         );
  HS65_GS_AND2X4 U954 ( .A(\mul_a1/fa1_s2_r[14] ), .B(\mul_a1/fa1_c1_r[13] ), 
        .Z(n907) );
  HS65_GSS_XOR2X3 U955 ( .A(\mul_a1/fa1_s1_r[15] ), .B(\mul_a1/fa1_s0_r[15] ), 
        .Z(n910) );
  HS65_GSS_XOR2X3 U956 ( .A(\mul_a1/fa1_s2_r[15] ), .B(\mul_a1/fa1_c1_r[14] ), 
        .Z(n909) );
  HS65_GS_AND2X4 U957 ( .A(\mul_a1/fa1_s1_r[14] ), .B(\mul_a1/fa1_s0_r[14] ), 
        .Z(n908) );
  HS65_GSS_XOR2X3 U958 ( .A(\mul_a1/fa1_s2_r[14] ), .B(\mul_a1/fa1_c1_r[13] ), 
        .Z(n865) );
  HS65_GSS_XOR2X3 U959 ( .A(\mul_a1/fa1_s1_r[14] ), .B(\mul_a1/fa1_s0_r[14] ), 
        .Z(n864) );
  HS65_GS_AND2X4 U960 ( .A(\mul_a1/fa1_s1_r[13] ), .B(\mul_a1/fa1_s0_r[13] ), 
        .Z(n863) );
  HS65_GS_IVX2 U961 ( .A(n902), .Z(n904) );
  HS65_GS_AND2X4 U962 ( .A(\mul_a1/fa1_s0_r[12] ), .B(\mul_a1/fa1_s1_r[12] ), 
        .Z(n867) );
  HS65_GSS_XOR2X3 U963 ( .A(\mul_a1/fa1_s1_r[13] ), .B(\mul_a1/fa1_s0_r[13] ), 
        .Z(n866) );
  HS65_GS_FA1X4 U964 ( .A0(n865), .B0(n864), .CI(n863), .CO(n905), .S0(n901)
         );
  HS65_GS_AND2X4 U965 ( .A(n900), .B(n901), .Z(n1771) );
  HS65_GSS_XOR2X3 U966 ( .A(\mul_a1/fa1_s0_r[11] ), .B(\mul_a1/fa1_s1_r[11] ), 
        .Z(n873) );
  HS65_GS_AND2X4 U967 ( .A(\mul_a1/fa1_s0_r[10] ), .B(\mul_a1/fa1_s1_r[10] ), 
        .Z(n872) );
  HS65_GSS_XOR2X3 U968 ( .A(\mul_a1/fa1_s0_r[12] ), .B(\mul_a1/fa1_s1_r[12] ), 
        .Z(n869) );
  HS65_GS_AND2X4 U969 ( .A(\mul_a1/fa1_s0_r[11] ), .B(\mul_a1/fa1_s1_r[11] ), 
        .Z(n868) );
  HS65_GS_AND2X4 U970 ( .A(n870), .B(n871), .Z(n895) );
  HS65_GS_FA1X4 U971 ( .A0(n867), .B0(\mul_a1/fa1_c1_r[12] ), .CI(n866), .CO(
        n900), .S0(n896) );
  HS65_GS_FA1X4 U972 ( .A0(\mul_a1/fa1_c1_r[11] ), .B0(n869), .CI(n868), .CO(
        n897), .S0(n871) );
  HS65_GSS_XOR2X3 U973 ( .A(n896), .B(n897), .Z(n894) );
  HS65_GSS_XOR2X3 U974 ( .A(n871), .B(n870), .Z(n892) );
  HS65_GSS_XOR2X3 U975 ( .A(\mul_a1/fa1_s0_r[10] ), .B(\mul_a1/fa1_s1_r[10] ), 
        .Z(n879) );
  HS65_GS_AND2X4 U976 ( .A(\mul_a1/fa1_s0_r[9] ), .B(\mul_a1/fa1_s1_r[9] ), 
        .Z(n878) );
  HS65_GS_FA1X4 U977 ( .A0(\mul_a1/fa1_c1_r[10] ), .B0(n873), .CI(n872), .CO(
        n870), .S0(n885) );
  HS65_GS_AND2X4 U978 ( .A(n884), .B(n885), .Z(n891) );
  HS65_GS_NAND2X2 U979 ( .A(\mul_a1/fa1_s0_r[7] ), .B(\mul_a1/fa1_s1_r[7] ), 
        .Z(n875) );
  HS65_GSS_XNOR2X3 U980 ( .A(\mul_a1/fa1_s1_r[8] ), .B(\mul_a1/fa1_s0_r[8] ), 
        .Z(n874) );
  HS65_GS_NOR2X2 U981 ( .A(n875), .B(n874), .Z(n877) );
  HS65_GS_AND2X4 U982 ( .A(\mul_a1/fa1_s1_r[8] ), .B(\mul_a1/fa1_s0_r[8] ), 
        .Z(n881) );
  HS65_GSS_XOR2X3 U983 ( .A(\mul_a1/fa1_s0_r[9] ), .B(\mul_a1/fa1_s1_r[9] ), 
        .Z(n880) );
  HS65_GS_NAND2X2 U984 ( .A(n877), .B(n876), .Z(n889) );
  HS65_GS_FA1X4 U985 ( .A0(\mul_a1/fa1_c1_r[9] ), .B0(n879), .CI(n878), .CO(
        n884), .S0(n883) );
  HS65_GS_IVX2 U986 ( .A(n883), .Z(n888) );
  HS65_GS_FA1X4 U987 ( .A0(n881), .B0(n880), .CI(\mul_a1/fa1_c1_r[8] ), .CO(
        n882), .S0(n876) );
  HS65_GS_NAND2X2 U988 ( .A(n883), .B(n882), .Z(n887) );
  HS65_GSS_XNOR2X3 U989 ( .A(n885), .B(n884), .Z(n886) );
  HS65_GS_CBI4I6X2 U990 ( .A(n889), .B(n888), .C(n887), .D(n886), .Z(n890) );
  HS65_GS_PAO2X4 U991 ( .A(n892), .B(n891), .P(n890), .Z(n893) );
  HS65_GS_PAOI2X1 U992 ( .A(n895), .B(n894), .P(n893), .Z(n899) );
  HS65_GS_AND2X4 U993 ( .A(n897), .B(n896), .Z(n898) );
  HS65_GS_NOR2AX3 U994 ( .A(n899), .B(n898), .Z(n1766) );
  HS65_GSS_XOR2X3 U995 ( .A(n901), .B(n900), .Z(n1767) );
  HS65_GS_NOR2X2 U996 ( .A(n1767), .B(n1766), .Z(n1765) );
  HS65_GS_NOR2X2 U997 ( .A(n1766), .B(n1765), .Z(n903) );
  HS65_GSS_XNOR2X3 U998 ( .A(n903), .B(n902), .Z(n1770) );
  HS65_GS_NOR2X2 U999 ( .A(n1771), .B(n1770), .Z(n1769) );
  HS65_GS_NOR2X2 U1000 ( .A(n904), .B(n1769), .Z(n912) );
  HS65_GS_FA1X4 U1001 ( .A0(n907), .B0(n906), .CI(n905), .CO(n911), .S0(n902)
         );
  HS65_GS_NOR2X2 U1002 ( .A(n912), .B(n911), .Z(n913) );
  HS65_GS_AND2X4 U1003 ( .A(\mul_a1/fa1_s2_r[15] ), .B(\mul_a1/fa1_c1_r[14] ), 
        .Z(n916) );
  HS65_GS_FA1X4 U1004 ( .A0(n910), .B0(n909), .CI(n908), .CO(n915), .S0(n906)
         );
  HS65_GSS_XOR2X3 U1005 ( .A(\mul_a1/fa1_s1_r[16] ), .B(\mul_a1/fa1_s0_r[16] ), 
        .Z(n919) );
  HS65_GSS_XOR2X3 U1006 ( .A(\mul_a1/fa1_s2_r[16] ), .B(\mul_a1/fa1_c1_r[15] ), 
        .Z(n918) );
  HS65_GS_AND2X4 U1007 ( .A(\mul_a1/fa1_s1_r[15] ), .B(\mul_a1/fa1_s0_r[15] ), 
        .Z(n917) );
  HS65_GSS_XNOR2X3 U1008 ( .A(n912), .B(n911), .Z(n1774) );
  HS65_GS_NOR2X2 U1009 ( .A(n1775), .B(n1774), .Z(n1773) );
  HS65_GS_NOR2X2 U1010 ( .A(n913), .B(n1773), .Z(n921) );
  HS65_GS_FA1X4 U1011 ( .A0(n916), .B0(n915), .CI(n914), .CO(n920), .S0(n1775)
         );
  HS65_GS_NOR2X2 U1012 ( .A(n921), .B(n920), .Z(n922) );
  HS65_GS_AND2X4 U1013 ( .A(\mul_a1/fa1_s2_r[16] ), .B(\mul_a1/fa1_c1_r[15] ), 
        .Z(n925) );
  HS65_GS_FA1X4 U1014 ( .A0(n919), .B0(n918), .CI(n917), .CO(n924), .S0(n914)
         );
  HS65_GSS_XOR2X3 U1015 ( .A(\mul_a1/fa1_s1_r[17] ), .B(\mul_a1/fa1_s0_r[17] ), 
        .Z(n928) );
  HS65_GSS_XOR2X3 U1016 ( .A(\mul_a1/fa1_s2_r[17] ), .B(\mul_a1/fa1_c1_r[16] ), 
        .Z(n927) );
  HS65_GS_AND2X4 U1017 ( .A(\mul_a1/fa1_s1_r[16] ), .B(\mul_a1/fa1_s0_r[16] ), 
        .Z(n926) );
  HS65_GSS_XNOR2X3 U1018 ( .A(n921), .B(n920), .Z(n1778) );
  HS65_GS_NOR2X2 U1019 ( .A(n1779), .B(n1778), .Z(n1777) );
  HS65_GS_NOR2X2 U1020 ( .A(n922), .B(n1777), .Z(n929) );
  HS65_GS_FA1X4 U1021 ( .A0(n925), .B0(n924), .CI(n923), .CO(n930), .S0(n1779)
         );
  HS65_GS_NOR2X2 U1022 ( .A(n929), .B(n930), .Z(n931) );
  HS65_GS_AND2X4 U1023 ( .A(\mul_a1/fa1_s2_r[17] ), .B(\mul_a1/fa1_c1_r[16] ), 
        .Z(n934) );
  HS65_GS_FA1X4 U1024 ( .A0(n928), .B0(n927), .CI(n926), .CO(n933), .S0(n923)
         );
  HS65_GSS_XOR2X3 U1025 ( .A(\mul_a1/fa1_s1_r[18] ), .B(\mul_a1/fa1_s0_r[18] ), 
        .Z(n937) );
  HS65_GSS_XOR2X3 U1026 ( .A(\mul_a1/fa1_s2_r[18] ), .B(\mul_a1/fa1_c1_r[17] ), 
        .Z(n936) );
  HS65_GS_AND2X4 U1027 ( .A(\mul_a1/fa1_s1_r[17] ), .B(\mul_a1/fa1_s0_r[17] ), 
        .Z(n935) );
  HS65_GSS_XNOR2X3 U1028 ( .A(n930), .B(n929), .Z(n1782) );
  HS65_GS_NOR2X2 U1029 ( .A(n1783), .B(n1782), .Z(n1781) );
  HS65_GS_NOR2X2 U1030 ( .A(n931), .B(n1781), .Z(n1653) );
  HS65_GS_FA1X4 U1031 ( .A0(n934), .B0(n933), .CI(n932), .CO(n1654), .S0(n1783) );
  HS65_GS_AND2X4 U1032 ( .A(\mul_a1/fa1_s2_r[18] ), .B(\mul_a1/fa1_c1_r[17] ), 
        .Z(n943) );
  HS65_GS_FA1X4 U1033 ( .A0(n937), .B0(n936), .CI(n935), .CO(n942), .S0(n932)
         );
  HS65_GS_FA1X4 U1034 ( .A0(n940), .B0(n939), .CI(n938), .CO(n861), .S0(n941)
         );
  HS65_GS_PAO2X4 U1035 ( .A(n1653), .B(n1654), .P(n1658), .Z(n1648) );
  HS65_GS_FA1X4 U1036 ( .A0(n943), .B0(n942), .CI(n941), .CO(n1649), .S0(n1658) );
  HS65_GS_PAO2X4 U1037 ( .A(n1652), .B(n1648), .P(n1649), .Z(n1644) );
  HS65_GS_FA1X4 U1038 ( .A0(n946), .B0(n945), .CI(n944), .CO(n1641), .S0(n1643) );
  HS65_GS_AND2X4 U1039 ( .A(\mul_a1/fa1_s2_r[21] ), .B(\mul_a1/fa1_c1_r[20] ), 
        .Z(n955) );
  HS65_GS_FA1X4 U1040 ( .A0(n949), .B0(n948), .CI(n947), .CO(n954), .S0(n944)
         );
  HS65_GS_FA1X4 U1041 ( .A0(n952), .B0(n951), .CI(n950), .CO(n957), .S0(n953)
         );
  HS65_GS_FA1X4 U1042 ( .A0(n955), .B0(n954), .CI(n953), .CO(n1636), .S0(n1639) );
  HS65_GS_FA1X4 U1043 ( .A0(n958), .B0(n957), .CI(n956), .CO(n1633), .S0(n1635) );
  HS65_GS_AND2X4 U1044 ( .A(\mul_a1/fa1_s2_r[23] ), .B(\mul_a1/fa1_c1_r[22] ), 
        .Z(n967) );
  HS65_GS_FA1X4 U1045 ( .A0(n961), .B0(n960), .CI(n959), .CO(n966), .S0(n956)
         );
  HS65_GS_FA1X4 U1046 ( .A0(n964), .B0(n963), .CI(n962), .CO(n969), .S0(n965)
         );
  HS65_GS_FA1X4 U1047 ( .A0(n967), .B0(n966), .CI(n965), .CO(n1628), .S0(n1631) );
  HS65_GS_FA1X4 U1048 ( .A0(n970), .B0(n969), .CI(n968), .CO(n1625), .S0(n1627) );
  HS65_GS_FA1X4 U1049 ( .A0(n973), .B0(n972), .CI(n971), .CO(n1621), .S0(n1623) );
  HS65_GS_FA1X4 U1050 ( .A0(n976), .B0(n975), .CI(n974), .CO(n1598), .S0(n1619) );
  HS65_GS_AND2X4 U1051 ( .A(\mul_a1/fa1_s2_r[27] ), .B(\mul_a1/fa1_c1_r[26] ), 
        .Z(n985) );
  HS65_GS_FA1X4 U1052 ( .A0(n979), .B0(n978), .CI(n977), .CO(n984), .S0(n974)
         );
  HS65_GS_FA1X4 U1053 ( .A0(n982), .B0(n981), .CI(n980), .CO(n987), .S0(n983)
         );
  HS65_GS_FA1X4 U1054 ( .A0(n985), .B0(n984), .CI(n983), .CO(n1603), .S0(n1596) );
  HS65_GS_FA1X4 U1055 ( .A0(n988), .B0(n987), .CI(n986), .CO(n1610), .S0(n1602) );
  HS65_GS_FA1X4 U1056 ( .A0(n991), .B0(n990), .CI(n989), .CO(n1607), .S0(n1608) );
  HS65_GS_AND2X4 U1057 ( .A(\mul_a1/fa1_s2_r[30] ), .B(\mul_a1/fa1_c1_r[29] ), 
        .Z(n1000) );
  HS65_GS_FA1X4 U1058 ( .A0(n994), .B0(n993), .CI(n992), .CO(n1001), .S0(n999)
         );
  HS65_GS_FA1X4 U1059 ( .A0(n997), .B0(n996), .CI(n995), .CO(n998), .S0(n989)
         );
  HS65_GS_FA1X4 U1060 ( .A0(n1000), .B0(n999), .CI(n998), .CO(n1599), .S0(
        n1605) );
  HS65_GS_FA1X4 U1061 ( .A0(n1003), .B0(n1002), .CI(n1001), .CO(n1012), .S0(
        n1601) );
  HS65_GS_FA1X4 U1062 ( .A0(n1006), .B0(n1005), .CI(n1004), .CO(n1010), .S0(
        n1002) );
  HS65_GS_NAND2X2 U1063 ( .A(\mul_a1/fa1_s2_r[32] ), .B(\mul_a1/fa1_c1_r[31] ), 
        .Z(n1009) );
  HS65_GSS_XOR3X2 U1064 ( .A(\mul_a1/fa1_s0_r[33] ), .B(\mul_a1/fa1_s2_r[33] ), 
        .C(n1007), .Z(n1008) );
  HS65_GSS_XOR3X2 U1065 ( .A(n1010), .B(n1009), .C(n1008), .Z(n1011) );
  HS65_GSS_XOR3X2 U1066 ( .A(n1013), .B(n1012), .C(n1011), .Z(n1014) );
  HS65_GSS_XOR3X2 U1067 ( .A(\mul_a1/fa1_s1_r[33] ), .B(\mul_a1/fa1_c1_r[32] ), 
        .C(n1014), .Z(\mul_a1/result_sat[15] ) );
  HS65_GS_IVX2 U1068 ( .A(x_reg2[14]), .Z(n1496) );
  HS65_GS_IVX2 U1069 ( .A(x_reg2[13]), .Z(n1498) );
  HS65_GS_IVX2 U1070 ( .A(x_reg2[12]), .Z(n1500) );
  HS65_GS_IVX2 U1071 ( .A(x_reg2[11]), .Z(n1502) );
  HS65_GS_IVX2 U1072 ( .A(x_reg2[10]), .Z(n1504) );
  HS65_GS_IVX2 U1073 ( .A(x_reg2[9]), .Z(n1506) );
  HS65_GS_IVX2 U1074 ( .A(x_reg2[8]), .Z(n1508) );
  HS65_GS_IVX2 U1075 ( .A(x_reg2[7]), .Z(n1510) );
  HS65_GS_IVX2 U1076 ( .A(x_reg2[6]), .Z(n1512) );
  HS65_GS_IVX2 U1077 ( .A(x_reg2[5]), .Z(n1514) );
  HS65_GS_IVX2 U1078 ( .A(x_reg2[4]), .Z(n1516) );
  HS65_GS_IVX2 U1079 ( .A(x_reg2[3]), .Z(n1518) );
  HS65_GS_IVX2 U1080 ( .A(x_reg2[2]), .Z(n1751) );
  HS65_GS_IVX2 U1081 ( .A(x_reg2[1]), .Z(n1742) );
  HS65_GS_IVX2 U1082 ( .A(x_reg2[0]), .Z(n1741) );
  HS65_GS_NOR2X3 U1083 ( .A(\DP_OP_371J1_181_1383/n79 ), .B(n1449), .Z(n1812)
         );
  HS65_GS_MUX21I1X3 U1084 ( .D0(n1753), .D1(data_out[0]), .S0(n1440), .Z(n1916) );
  HS65_GS_IVX2 U1085 ( .A(x_z1[14]), .Z(n1436) );
  HS65_GS_IVX2 U1086 ( .A(x_z1[13]), .Z(n1435) );
  HS65_GS_IVX2 U1087 ( .A(x_z1[12]), .Z(n1433) );
  HS65_GS_IVX2 U1088 ( .A(x_z1[11]), .Z(n1431) );
  HS65_GS_IVX2 U1089 ( .A(x_z1[10]), .Z(n1430) );
  HS65_GS_IVX2 U1090 ( .A(x_z1[9]), .Z(n1427) );
  HS65_GS_IVX2 U1091 ( .A(x_z1[8]), .Z(n1426) );
  HS65_GS_IVX2 U1092 ( .A(x_z1[7]), .Z(n1424) );
  HS65_GS_IVX2 U1093 ( .A(x_z1[6]), .Z(n1422) );
  HS65_GS_IVX2 U1094 ( .A(x_z1[5]), .Z(n1420) );
  HS65_GS_IVX2 U1095 ( .A(x_z1[4]), .Z(n1417) );
  HS65_GS_IVX2 U1096 ( .A(x_z1[3]), .Z(n1415) );
  HS65_GS_IVX2 U1097 ( .A(x_z1[2]), .Z(n1413) );
  HS65_GS_IVX2 U1098 ( .A(x_z1[1]), .Z(n1412) );
  HS65_GS_IVX2 U1099 ( .A(x_z1[0]), .Z(n1410) );
  HS65_GS_NOR2X2 U1100 ( .A(x_z1[15]), .B(n1016), .Z(n1015) );
  HS65_GSS_XNOR2X3 U1101 ( .A(n1015), .B(n1438), .Z(\mul_b0/fa1_s0[30] ) );
  HS65_GSS_XNOR2X3 U1102 ( .A(x_z1[15]), .B(n1016), .Z(n1119) );
  HS65_GSS_XNOR2X3 U1103 ( .A(n1119), .B(n1438), .Z(\mul_b0/fa1_s0[20] ) );
  HS65_GSS_XOR2X3 U1104 ( .A(n1310), .B(y_z2[1]), .Z(\mul_a2/fa1_s0[3] ) );
  HS65_GS_NOR2X2 U1105 ( .A(\DP_OP_371J1_181_1383/n79 ), .B(n1492), .Z(n1519)
         );
  HS65_GSS_XNOR2X3 U1106 ( .A(n1519), .B(n1494), .Z(\mul_b2/fa1_s1[28] ) );
  HS65_GS_BFX4 U1107 ( .A(n1821), .Z(n1437) );
  HS65_GS_MUXI21X2 U1108 ( .D0(n1701), .D1(n1753), .S0(n1437), .Z(n1917) );
  HS65_GS_IVX2 U1109 ( .A(x_z2[0]), .Z(n1411) );
  HS65_GSS_XNOR2X3 U1110 ( .A(n1583), .B(n1749), .Z(\mul_b1/fa1_s2[26] ) );
  HS65_GS_HA1X4 U1111 ( .A0(n1749), .B0(n1017), .CO(n1116), .S0(n1584) );
  HS65_GSS_XNOR2X3 U1112 ( .A(n1584), .B(n1432), .Z(\mul_b1/fa1_s2[25] ) );
  HS65_GS_HA1X4 U1113 ( .A0(n1432), .B0(n1018), .CO(n1017), .S0(n1585) );
  HS65_GSS_XNOR2X3 U1114 ( .A(n1585), .B(n1429), .Z(\mul_b1/fa1_s2[24] ) );
  HS65_GS_HA1X4 U1115 ( .A0(n1429), .B0(n1019), .CO(n1018), .S0(n1586) );
  HS65_GSS_XNOR2X3 U1116 ( .A(n1586), .B(n1428), .Z(\mul_b1/fa1_s2[23] ) );
  HS65_GS_HA1X4 U1117 ( .A0(n1428), .B0(n1020), .CO(n1019), .S0(n1587) );
  HS65_GSS_XNOR2X3 U1118 ( .A(n1587), .B(n1425), .Z(\mul_b1/fa1_s2[22] ) );
  HS65_GS_HA1X4 U1119 ( .A0(n1425), .B0(n1021), .CO(n1020), .S0(n1588) );
  HS65_GSS_XNOR2X3 U1120 ( .A(n1588), .B(n1423), .Z(\mul_b1/fa1_s2[21] ) );
  HS65_GS_HA1X4 U1121 ( .A0(n1423), .B0(n1022), .CO(n1021), .S0(n1589) );
  HS65_GSS_XNOR2X3 U1122 ( .A(n1589), .B(n1421), .Z(\mul_b1/fa1_s2[20] ) );
  HS65_GS_HA1X4 U1123 ( .A0(n1421), .B0(n1023), .CO(n1022), .S0(n1590) );
  HS65_GSS_XNOR2X3 U1124 ( .A(n1590), .B(n1419), .Z(\mul_b1/fa1_s2[19] ) );
  HS65_GS_HA1X4 U1125 ( .A0(n1419), .B0(n1024), .CO(n1023), .S0(n1591) );
  HS65_GSS_XNOR2X3 U1126 ( .A(n1591), .B(n1418), .Z(\mul_b1/fa1_s2[18] ) );
  HS65_GS_HA1X4 U1127 ( .A0(n1418), .B0(n1025), .CO(n1024), .S0(n1592) );
  HS65_GSS_XNOR2X3 U1128 ( .A(n1592), .B(n1416), .Z(\mul_b1/fa1_s2[17] ) );
  HS65_GS_HA1X4 U1129 ( .A0(n1416), .B0(n1026), .CO(n1025), .S0(n1593) );
  HS65_GSS_XNOR2X3 U1130 ( .A(n1593), .B(n1414), .Z(\mul_b1/fa1_s2[16] ) );
  HS65_GS_HA1X4 U1131 ( .A0(n1414), .B0(n1027), .CO(n1026), .S0(n1594) );
  HS65_GSS_XNOR2X3 U1132 ( .A(n1594), .B(n1752), .Z(\mul_b1/fa1_s2[15] ) );
  HS65_GS_HA1X4 U1133 ( .A0(n1752), .B0(n1411), .CO(n1027), .S0(n1595) );
  HS65_GSS_XNOR2X3 U1134 ( .A(n1595), .B(n1411), .Z(\mul_b1/fa1_s2[14] ) );
  HS65_GS_FA1X4 U1135 ( .A0(n1030), .B0(n1029), .CI(n1028), .CO(n1036), .S0(
        n1050) );
  HS65_GS_FA1X4 U1136 ( .A0(n1033), .B0(n1032), .CI(n1031), .CO(n1042), .S0(
        n1049) );
  HS65_GS_FA1X4 U1137 ( .A0(n1036), .B0(n1035), .CI(n1034), .CO(n1032), .S0(
        n1046) );
  HS65_GS_FA1X4 U1138 ( .A0(n1039), .B0(n1038), .CI(n1037), .CO(n606), .S0(
        n1045) );
  HS65_GS_FA1X4 U1139 ( .A0(n1042), .B0(n1041), .CI(n1040), .CO(n1038), .S0(
        n1044) );
  HS65_GS_AND3X4 U1140 ( .A(n1046), .B(n1045), .C(n1044), .Z(n1043) );
  HS65_GS_IVX2 U1141 ( .A(\mul_b1/result_sat[15] ), .Z(n1047) );
  HS65_GS_AOI12X2 U1142 ( .A(n1049), .B(n1043), .C(n1047), .Z(n1796) );
  HS65_GS_IVX2 U1143 ( .A(n1796), .Z(n1103) );
  HS65_GS_OR3X4 U1144 ( .A(n1046), .B(n1045), .C(n1044), .Z(n1048) );
  HS65_GS_OAI21X2 U1145 ( .A(n1049), .B(n1048), .C(n1047), .Z(n1797) );
  HS65_GS_IVX2 U1146 ( .A(n1797), .Z(n1102) );
  HS65_GS_AO12X4 U1147 ( .A(n1050), .B(n1103), .C(n1102), .Z(
        \mul_b1/result_sat[14] ) );
  HS65_GS_FA1X4 U1148 ( .A0(n1053), .B0(n1052), .CI(n1051), .CO(n1029), .S0(
        n1054) );
  HS65_GS_OA12X4 U1149 ( .A(n1102), .B(n1054), .C(n1103), .Z(
        \mul_b1/result_sat[13] ) );
  HS65_GS_FA1X4 U1150 ( .A0(n1057), .B0(n1056), .CI(n1055), .CO(n1052), .S0(
        n1058) );
  HS65_GS_AO12X4 U1151 ( .A(n1058), .B(n1103), .C(n1102), .Z(
        \mul_b1/result_sat[12] ) );
  HS65_GS_FA1X4 U1152 ( .A0(n1061), .B0(n1060), .CI(n1059), .CO(n1057), .S0(
        n1062) );
  HS65_GS_AO12X4 U1153 ( .A(n1062), .B(n1103), .C(n1102), .Z(
        \mul_b1/result_sat[11] ) );
  HS65_GS_FA1X4 U1154 ( .A0(n1065), .B0(n1064), .CI(n1063), .CO(n1061), .S0(
        n1066) );
  HS65_GS_OA12X4 U1155 ( .A(n1102), .B(n1066), .C(n1103), .Z(
        \mul_b1/result_sat[10] ) );
  HS65_GS_FA1X4 U1156 ( .A0(n1069), .B0(n1068), .CI(n1067), .CO(n1064), .S0(
        n1070) );
  HS65_GS_OA12X4 U1157 ( .A(n1102), .B(n1070), .C(n1103), .Z(
        \mul_b1/result_sat[9] ) );
  HS65_GS_FA1X4 U1158 ( .A0(n1073), .B0(n1072), .CI(n1071), .CO(n1068), .S0(
        n1074) );
  HS65_GS_AO12X4 U1159 ( .A(n1074), .B(n1103), .C(n1102), .Z(
        \mul_b1/result_sat[8] ) );
  HS65_GS_FA1X4 U1160 ( .A0(n1077), .B0(n1076), .CI(n1075), .CO(n1073), .S0(
        n1078) );
  HS65_GS_AO12X4 U1161 ( .A(n1078), .B(n1103), .C(n1102), .Z(
        \mul_b1/result_sat[7] ) );
  HS65_GS_FA1X4 U1162 ( .A0(n1081), .B0(n1080), .CI(n1079), .CO(n1076), .S0(
        n1082) );
  HS65_GS_OA12X4 U1163 ( .A(n1102), .B(n1082), .C(n1103), .Z(
        \mul_b1/result_sat[6] ) );
  HS65_GS_FA1X4 U1164 ( .A0(n1085), .B0(n1084), .CI(n1083), .CO(n1080), .S0(
        n1086) );
  HS65_GS_AO12X4 U1165 ( .A(n1086), .B(n1103), .C(n1102), .Z(
        \mul_b1/result_sat[5] ) );
  HS65_GS_FA1X4 U1166 ( .A0(n1089), .B0(n1088), .CI(n1087), .CO(n1084), .S0(
        n1090) );
  HS65_GS_AO12X4 U1167 ( .A(n1090), .B(n1103), .C(n1102), .Z(
        \mul_b1/result_sat[4] ) );
  HS65_GS_FA1X4 U1168 ( .A0(n1093), .B0(n1092), .CI(n1091), .CO(n1088), .S0(
        n1094) );
  HS65_GS_OA12X4 U1169 ( .A(n1102), .B(n1094), .C(n1103), .Z(
        \mul_b1/result_sat[3] ) );
  HS65_GS_FA1X4 U1170 ( .A0(n1097), .B0(n1096), .CI(n1095), .CO(n1093), .S0(
        n1098) );
  HS65_GS_AO12X4 U1171 ( .A(n1098), .B(n1103), .C(n1102), .Z(
        \mul_b1/result_sat[2] ) );
  HS65_GS_FA1X4 U1172 ( .A0(n1101), .B0(n1100), .CI(n1099), .CO(n1097), .S0(
        n1104) );
  HS65_GS_AO12X4 U1173 ( .A(n1104), .B(n1103), .C(n1102), .Z(
        \mul_b1/result_sat[1] ) );
  HS65_GS_HA1X4 U1174 ( .A0(n1436), .B0(n1105), .CO(n1016), .S0(n1120) );
  HS65_GSS_XNOR2X3 U1175 ( .A(n1120), .B(n1438), .Z(\mul_b0/fa1_s0[19] ) );
  HS65_GS_HA1X4 U1176 ( .A0(n1435), .B0(n1106), .CO(n1105), .S0(n1121) );
  HS65_GSS_XNOR2X3 U1177 ( .A(n1121), .B(n1438), .Z(\mul_b0/fa1_s0[18] ) );
  HS65_GS_HA1X4 U1178 ( .A0(n1433), .B0(n1107), .CO(n1106), .S0(n1122) );
  HS65_GSS_XNOR2X3 U1179 ( .A(n1122), .B(n1438), .Z(\mul_b0/fa1_s0[17] ) );
  HS65_GS_HA1X4 U1180 ( .A0(n1431), .B0(n1108), .CO(n1107), .S0(n1123) );
  HS65_GSS_XNOR2X3 U1181 ( .A(n1123), .B(n1438), .Z(\mul_b0/fa1_s0[16] ) );
  HS65_GS_HA1X4 U1182 ( .A0(n1430), .B0(n1109), .CO(n1108), .S0(n1124) );
  HS65_GSS_XNOR2X3 U1183 ( .A(n1124), .B(n1438), .Z(\mul_b0/fa1_s0[15] ) );
  HS65_GS_HA1X4 U1184 ( .A0(n1427), .B0(n1110), .CO(n1109), .S0(n1125) );
  HS65_GSS_XNOR2X3 U1185 ( .A(n1125), .B(n1436), .Z(\mul_b0/fa1_s0[14] ) );
  HS65_GS_HA1X4 U1186 ( .A0(n1426), .B0(n1111), .CO(n1110), .S0(n1126) );
  HS65_GSS_XNOR2X3 U1187 ( .A(n1126), .B(n1435), .Z(\mul_b0/fa1_s0[13] ) );
  HS65_GS_HA1X4 U1188 ( .A0(n1424), .B0(n1112), .CO(n1111), .S0(n1127) );
  HS65_GSS_XNOR2X3 U1189 ( .A(n1127), .B(n1433), .Z(\mul_b0/fa1_s0[12] ) );
  HS65_GS_HA1X4 U1190 ( .A0(n1422), .B0(n1113), .CO(n1112), .S0(n1128) );
  HS65_GSS_XNOR2X3 U1191 ( .A(n1128), .B(n1431), .Z(\mul_b0/fa1_s0[11] ) );
  HS65_GS_HA1X4 U1192 ( .A0(n1420), .B0(n1114), .CO(n1113), .S0(n1129) );
  HS65_GSS_XNOR2X3 U1193 ( .A(n1129), .B(n1430), .Z(\mul_b0/fa1_s0[10] ) );
  HS65_GS_HA1X4 U1194 ( .A0(n1417), .B0(n1115), .CO(n1114), .S0(n1130) );
  HS65_GSS_XNOR2X3 U1195 ( .A(n1130), .B(n1427), .Z(\mul_b0/fa1_s0[9] ) );
  HS65_GS_HA1X4 U1196 ( .A0(n1747), .B0(n1116), .CO(n1175), .S0(n1583) );
  HS65_GSS_XNOR2X3 U1197 ( .A(n1582), .B(n1747), .Z(\mul_b1/fa1_s2[27] ) );
  HS65_GS_HA1X4 U1198 ( .A0(n1415), .B0(n1117), .CO(n1115), .S0(n1131) );
  HS65_GSS_XNOR2X3 U1199 ( .A(n1131), .B(n1426), .Z(\mul_b0/fa1_s0[8] ) );
  HS65_GS_HA1X4 U1200 ( .A0(n1413), .B0(n1118), .CO(n1117), .S0(n1132) );
  HS65_GSS_XNOR2X3 U1201 ( .A(n1132), .B(n1424), .Z(\mul_b0/fa1_s0[7] ) );
  HS65_GS_HA1X4 U1202 ( .A0(n1412), .B0(n1410), .CO(n1118), .S0(n1133) );
  HS65_GSS_XNOR2X3 U1203 ( .A(n1133), .B(n1422), .Z(\mul_b0/fa1_s0[6] ) );
  HS65_GS_AND2X4 U1204 ( .A(n1119), .B(n1820), .Z(\mul_b0/fa1_c0[20] ) );
  HS65_GS_AND2X4 U1205 ( .A(n1120), .B(x_z1[15]), .Z(\mul_b0/fa1_c0[19] ) );
  HS65_GS_AND2X4 U1206 ( .A(n1121), .B(n1820), .Z(\mul_b0/fa1_c0[18] ) );
  HS65_GS_AND2X4 U1207 ( .A(n1122), .B(x_z1[15]), .Z(\mul_b0/fa1_c0[17] ) );
  HS65_GS_AND2X4 U1208 ( .A(n1123), .B(n1820), .Z(\mul_b0/fa1_c0[16] ) );
  HS65_GS_AND2X4 U1209 ( .A(n1124), .B(x_z1[15]), .Z(\mul_b0/fa1_c0[15] ) );
  HS65_GS_AND2X4 U1210 ( .A(n1125), .B(x_z1[14]), .Z(\mul_b0/fa1_c0[14] ) );
  HS65_GS_AND2X4 U1211 ( .A(n1126), .B(x_z1[13]), .Z(\mul_b0/fa1_c0[13] ) );
  HS65_GS_AND2X4 U1212 ( .A(n1127), .B(x_z1[12]), .Z(\mul_b0/fa1_c0[12] ) );
  HS65_GS_AND2X4 U1213 ( .A(n1128), .B(x_z1[11]), .Z(\mul_b0/fa1_c0[11] ) );
  HS65_GS_AND2X4 U1214 ( .A(n1129), .B(x_z1[10]), .Z(\mul_b0/fa1_c0[10] ) );
  HS65_GS_AND2X4 U1215 ( .A(n1130), .B(x_z1[9]), .Z(\mul_b0/fa1_c0[9] ) );
  HS65_GS_AND2X4 U1216 ( .A(x_z1[8]), .B(n1131), .Z(\mul_b0/fa1_c0[8] ) );
  HS65_GS_AND2X4 U1217 ( .A(n1132), .B(x_z1[7]), .Z(\mul_b0/fa1_c0[7] ) );
  HS65_GS_AND2X4 U1218 ( .A(x_z1[6]), .B(n1133), .Z(\mul_b0/fa1_c0[6] ) );
  HS65_GS_AND2X4 U1219 ( .A(x_z1[0]), .B(x_z1[5]), .Z(\mul_b0/fa1_c0[5] ) );
  HS65_GS_FA1X4 U1220 ( .A0(n1136), .B0(n1135), .CI(n1134), .CO(n619), .S0(
        n1137) );
  HS65_GS_AO12X4 U1221 ( .A(n1137), .B(n1167), .C(n1166), .Z(
        \mul_b0/result_sat[14] ) );
  HS65_GS_FA1X4 U1222 ( .A0(n1140), .B0(n1139), .CI(n1138), .CO(n1136), .S0(
        n1141) );
  HS65_GS_AO12X4 U1223 ( .A(n1141), .B(n1167), .C(n1166), .Z(
        \mul_b0/result_sat[13] ) );
  HS65_GS_FA1X4 U1224 ( .A0(n1144), .B0(n1143), .CI(n1142), .CO(n1138), .S0(
        n1145) );
  HS65_GS_OA12X4 U1225 ( .A(n1166), .B(n1145), .C(n1167), .Z(
        \mul_b0/result_sat[12] ) );
  HS65_GS_FA1X4 U1226 ( .A0(n1148), .B0(n1147), .CI(n1146), .CO(n632), .S0(
        n1149) );
  HS65_GS_AO12X4 U1227 ( .A(n1149), .B(n1167), .C(n1166), .Z(
        \mul_b0/result_sat[10] ) );
  HS65_GS_FA1X4 U1228 ( .A0(n1152), .B0(n1151), .CI(n1150), .CO(n1148), .S0(
        n1153) );
  HS65_GS_AO12X4 U1229 ( .A(n1153), .B(n1167), .C(n1166), .Z(
        \mul_b0/result_sat[9] ) );
  HS65_GS_FA1X4 U1230 ( .A0(n1156), .B0(n1155), .CI(n1154), .CO(n1152), .S0(
        n1157) );
  HS65_GS_AO12X4 U1231 ( .A(n1157), .B(n1167), .C(n1166), .Z(
        \mul_b0/result_sat[8] ) );
  HS65_GS_FA1X4 U1232 ( .A0(n1160), .B0(n1159), .CI(n1158), .CO(n1156), .S0(
        n1161) );
  HS65_GS_AO12X4 U1233 ( .A(n1161), .B(n1167), .C(n1166), .Z(
        \mul_b0/result_sat[7] ) );
  HS65_GS_FA1X4 U1234 ( .A0(n1164), .B0(n1163), .CI(n1162), .CO(n1158), .S0(
        n1165) );
  HS65_GS_OA12X4 U1235 ( .A(n1166), .B(n1165), .C(n1167), .Z(
        \mul_b0/result_sat[6] ) );
  HS65_GS_IVX2 U1236 ( .A(n1167), .Z(n1805) );
  HS65_GS_OAI21X2 U1237 ( .A(n1170), .B(n1169), .C(n1168), .Z(n1171) );
  HS65_GS_OAI21X2 U1238 ( .A(n1805), .B(n1171), .C(n1806), .Z(
        \mul_b0/result_sat[3] ) );
  HS65_GS_OAI21X2 U1239 ( .A(n1173), .B(n1172), .C(n1800), .Z(n1174) );
  HS65_GS_OAI21X2 U1240 ( .A(n1805), .B(n1174), .C(n1806), .Z(
        \mul_b0/result_sat[0] ) );
  HS65_GS_HA1X4 U1241 ( .A0(n1745), .B0(n1175), .CO(n1282), .S0(n1582) );
  HS65_GSS_XNOR2X3 U1242 ( .A(\DP_OP_331J1_157_5454/n87 ), .B(n1282), .Z(n1581) );
  HS65_GSS_XNOR2X3 U1243 ( .A(n1581), .B(n1745), .Z(\mul_b1/fa1_s2[28] ) );
  HS65_GS_HA1X4 U1244 ( .A0(n1432), .B0(n1176), .CO(n1748), .S0(n1186) );
  HS65_GSS_XOR3X2 U1245 ( .A(\DP_OP_331J1_157_5454/n87 ), .B(x_z2[14]), .C(
        n1186), .Z(\mul_b1/fa1_s0[16] ) );
  HS65_GS_HA1X4 U1246 ( .A0(n1429), .B0(n1177), .CO(n1176), .S0(n1189) );
  HS65_GSS_XOR3X2 U1247 ( .A(\DP_OP_331J1_157_5454/n87 ), .B(x_z2[13]), .C(
        n1189), .Z(\mul_b1/fa1_s0[15] ) );
  HS65_GS_HA1X4 U1248 ( .A0(n1428), .B0(n1178), .CO(n1177), .S0(n1192) );
  HS65_GSS_XOR3X2 U1249 ( .A(x_z2[12]), .B(x_z2[14]), .C(n1192), .Z(
        \mul_b1/fa1_s0[14] ) );
  HS65_GS_HA1X4 U1250 ( .A0(n1425), .B0(n1179), .CO(n1178), .S0(n1195) );
  HS65_GSS_XOR3X2 U1251 ( .A(x_z2[11]), .B(x_z2[13]), .C(n1195), .Z(
        \mul_b1/fa1_s0[13] ) );
  HS65_GS_HA1X4 U1252 ( .A0(n1423), .B0(n1180), .CO(n1179), .S0(n1198) );
  HS65_GSS_XOR3X2 U1253 ( .A(x_z2[10]), .B(x_z2[12]), .C(n1198), .Z(
        \mul_b1/fa1_s0[12] ) );
  HS65_GS_HA1X4 U1254 ( .A0(n1421), .B0(n1181), .CO(n1180), .S0(n1201) );
  HS65_GSS_XOR3X2 U1255 ( .A(x_z2[11]), .B(x_z2[9]), .C(n1201), .Z(
        \mul_b1/fa1_s0[11] ) );
  HS65_GS_HA1X4 U1256 ( .A0(n1419), .B0(n1182), .CO(n1181), .S0(n1204) );
  HS65_GSS_XOR3X2 U1257 ( .A(x_z2[10]), .B(x_z2[8]), .C(n1204), .Z(
        \mul_b1/fa1_s0[10] ) );
  HS65_GS_HA1X4 U1258 ( .A0(n1418), .B0(n1183), .CO(n1182), .S0(n1207) );
  HS65_GSS_XOR3X2 U1259 ( .A(x_z2[9]), .B(x_z2[7]), .C(n1207), .Z(
        \mul_b1/fa1_s0[9] ) );
  HS65_GS_HA1X4 U1260 ( .A0(n1416), .B0(n1184), .CO(n1183), .S0(n1210) );
  HS65_GSS_XOR3X2 U1261 ( .A(x_z2[8]), .B(x_z2[6]), .C(n1210), .Z(
        \mul_b1/fa1_s0[8] ) );
  HS65_GS_HA1X4 U1262 ( .A0(n1414), .B0(n1185), .CO(n1184), .S0(n1213) );
  HS65_GSS_XOR3X2 U1263 ( .A(x_z2[7]), .B(x_z2[5]), .C(n1213), .Z(
        \mul_b1/fa1_s0[7] ) );
  HS65_GS_HA1X4 U1264 ( .A0(n1752), .B0(n1411), .CO(n1185), .S0(n1216) );
  HS65_GSS_XOR3X2 U1265 ( .A(x_z2[6]), .B(x_z2[4]), .C(n1216), .Z(
        \mul_b1/fa1_s0[6] ) );
  HS65_GSS_XOR3X2 U1266 ( .A(x_z2[5]), .B(x_z2[3]), .C(x_z2[0]), .Z(
        \mul_b1/fa1_s0[5] ) );
  HS65_GS_IVX2 U1267 ( .A(n1186), .Z(n1188) );
  HS65_GS_OAI21X2 U1268 ( .A(\DP_OP_331J1_157_5454/n87 ), .B(n1186), .C(
        x_z2[14]), .Z(n1187) );
  HS65_GS_OAI21X2 U1269 ( .A(n1439), .B(n1188), .C(n1187), .Z(
        \mul_b1/fa1_c0[16] ) );
  HS65_GS_IVX2 U1270 ( .A(n1189), .Z(n1191) );
  HS65_GS_OAI21X2 U1271 ( .A(\DP_OP_331J1_157_5454/n87 ), .B(n1189), .C(
        x_z2[13]), .Z(n1190) );
  HS65_GS_OAI21X2 U1272 ( .A(n1439), .B(n1191), .C(n1190), .Z(
        \mul_b1/fa1_c0[15] ) );
  HS65_GS_IVX2 U1273 ( .A(n1192), .Z(n1194) );
  HS65_GS_OAI21X2 U1274 ( .A(x_z2[14]), .B(n1192), .C(x_z2[12]), .Z(n1193) );
  HS65_GS_OAI21X2 U1275 ( .A(n1745), .B(n1194), .C(n1193), .Z(
        \mul_b1/fa1_c0[14] ) );
  HS65_GS_IVX2 U1276 ( .A(n1195), .Z(n1197) );
  HS65_GS_OAI21X2 U1277 ( .A(x_z2[13]), .B(n1195), .C(x_z2[11]), .Z(n1196) );
  HS65_GS_OAI21X2 U1278 ( .A(n1747), .B(n1197), .C(n1196), .Z(
        \mul_b1/fa1_c0[13] ) );
  HS65_GS_IVX2 U1279 ( .A(n1198), .Z(n1200) );
  HS65_GS_OAI21X2 U1280 ( .A(x_z2[12]), .B(n1198), .C(x_z2[10]), .Z(n1199) );
  HS65_GS_OAI21X2 U1281 ( .A(n1749), .B(n1200), .C(n1199), .Z(
        \mul_b1/fa1_c0[12] ) );
  HS65_GS_IVX2 U1282 ( .A(n1201), .Z(n1203) );
  HS65_GS_OAI21X2 U1283 ( .A(x_z2[11]), .B(n1201), .C(x_z2[9]), .Z(n1202) );
  HS65_GS_OAI21X2 U1284 ( .A(n1432), .B(n1203), .C(n1202), .Z(
        \mul_b1/fa1_c0[11] ) );
  HS65_GS_IVX2 U1285 ( .A(n1204), .Z(n1206) );
  HS65_GS_OAI21X2 U1286 ( .A(x_z2[10]), .B(n1204), .C(x_z2[8]), .Z(n1205) );
  HS65_GS_OAI21X2 U1287 ( .A(n1429), .B(n1206), .C(n1205), .Z(
        \mul_b1/fa1_c0[10] ) );
  HS65_GS_IVX2 U1288 ( .A(n1207), .Z(n1209) );
  HS65_GS_OAI21X2 U1289 ( .A(x_z2[9]), .B(n1207), .C(x_z2[7]), .Z(n1208) );
  HS65_GS_OAI21X2 U1290 ( .A(n1428), .B(n1209), .C(n1208), .Z(
        \mul_b1/fa1_c0[9] ) );
  HS65_GS_IVX2 U1291 ( .A(n1210), .Z(n1212) );
  HS65_GS_OAI21X2 U1292 ( .A(x_z2[8]), .B(n1210), .C(x_z2[6]), .Z(n1211) );
  HS65_GS_OAI21X2 U1293 ( .A(n1425), .B(n1212), .C(n1211), .Z(
        \mul_b1/fa1_c0[8] ) );
  HS65_GS_IVX2 U1294 ( .A(n1213), .Z(n1215) );
  HS65_GS_OAI21X2 U1295 ( .A(x_z2[7]), .B(n1213), .C(x_z2[5]), .Z(n1214) );
  HS65_GS_OAI21X2 U1296 ( .A(n1423), .B(n1215), .C(n1214), .Z(
        \mul_b1/fa1_c0[7] ) );
  HS65_GS_IVX2 U1297 ( .A(n1216), .Z(n1218) );
  HS65_GS_OAI21X2 U1298 ( .A(x_z2[6]), .B(n1216), .C(x_z2[4]), .Z(n1217) );
  HS65_GS_OAI21X2 U1299 ( .A(n1421), .B(n1218), .C(n1217), .Z(
        \mul_b1/fa1_c0[6] ) );
  HS65_GS_OAI21X2 U1300 ( .A(x_z2[5]), .B(x_z2[0]), .C(x_z2[3]), .Z(n1219) );
  HS65_GS_OAI21X2 U1301 ( .A(n1419), .B(n1411), .C(n1219), .Z(
        \mul_b1/fa1_c0[5] ) );
  HS65_GS_NOR2X2 U1302 ( .A(\DP_OP_331J1_157_5454/n87 ), .B(n1221), .Z(n1220)
         );
  HS65_GSS_XOR3X2 U1303 ( .A(n1220), .B(\DP_OP_331J1_157_5454/n87 ), .C(n1), 
        .Z(\mul_b1/fa1_s1[25] ) );
  HS65_GSS_XNOR2X3 U1304 ( .A(\DP_OP_331J1_157_5454/n87 ), .B(n1221), .Z(n1222) );
  HS65_GSS_XOR3X2 U1305 ( .A(n1), .B(x_z2[14]), .C(n1222), .Z(
        \mul_b1/fa1_s1[24] ) );
  HS65_GS_HA1X4 U1306 ( .A0(n1439), .B0(n1223), .CO(n1221), .S0(n1224) );
  HS65_GSS_XOR3X2 U1307 ( .A(n1), .B(x_z2[13]), .C(n1224), .Z(
        \mul_b1/fa1_s1[23] ) );
  HS65_GSS_XNOR2X3 U1308 ( .A(\DP_OP_331J1_157_5454/n87 ), .B(n1225), .Z(n1254) );
  HS65_GS_HA1X4 U1309 ( .A0(n1745), .B0(n1226), .CO(n1223), .S0(n1253) );
  HS65_GSS_XOR3X2 U1310 ( .A(x_z2[12]), .B(n1254), .C(n1253), .Z(
        \mul_b1/fa1_s1[22] ) );
  HS65_GS_HA1X4 U1311 ( .A0(n1439), .B0(n1227), .CO(n1225), .S0(n1256) );
  HS65_GS_HA1X4 U1312 ( .A0(n1747), .B0(n1228), .CO(n1226), .S0(n1255) );
  HS65_GSS_XOR3X2 U1313 ( .A(x_z2[11]), .B(n1256), .C(n1255), .Z(
        \mul_b1/fa1_s1[21] ) );
  HS65_GS_HA1X4 U1314 ( .A0(n1745), .B0(n1229), .CO(n1227), .S0(n1258) );
  HS65_GS_HA1X4 U1315 ( .A0(n1749), .B0(n1230), .CO(n1228), .S0(n1257) );
  HS65_GSS_XOR3X2 U1316 ( .A(x_z2[10]), .B(n1258), .C(n1257), .Z(
        \mul_b1/fa1_s1[20] ) );
  HS65_GS_HA1X4 U1317 ( .A0(n1432), .B0(n1231), .CO(n1230), .S0(n1260) );
  HS65_GS_HA1X4 U1318 ( .A0(n1747), .B0(n1232), .CO(n1229), .S0(n1259) );
  HS65_GSS_XOR3X2 U1319 ( .A(x_z2[9]), .B(n1260), .C(n1259), .Z(
        \mul_b1/fa1_s1[19] ) );
  HS65_GS_HA1X4 U1320 ( .A0(n1749), .B0(n1233), .CO(n1232), .S0(n1262) );
  HS65_GS_HA1X4 U1321 ( .A0(n1429), .B0(n1234), .CO(n1231), .S0(n1261) );
  HS65_GSS_XOR3X2 U1322 ( .A(x_z2[8]), .B(n1262), .C(n1261), .Z(
        \mul_b1/fa1_s1[18] ) );
  HS65_GS_HA1X4 U1323 ( .A0(n1432), .B0(n1235), .CO(n1233), .S0(n1264) );
  HS65_GS_HA1X4 U1324 ( .A0(n1428), .B0(n1236), .CO(n1234), .S0(n1263) );
  HS65_GSS_XOR3X2 U1325 ( .A(x_z2[7]), .B(n1264), .C(n1263), .Z(
        \mul_b1/fa1_s1[17] ) );
  HS65_GS_HA1X4 U1326 ( .A0(n1429), .B0(n1237), .CO(n1235), .S0(n1266) );
  HS65_GS_HA1X4 U1327 ( .A0(n1425), .B0(n1238), .CO(n1236), .S0(n1265) );
  HS65_GSS_XOR3X2 U1328 ( .A(x_z2[6]), .B(n1266), .C(n1265), .Z(
        \mul_b1/fa1_s1[16] ) );
  HS65_GS_HA1X4 U1329 ( .A0(n1428), .B0(n1239), .CO(n1237), .S0(n1268) );
  HS65_GS_HA1X4 U1330 ( .A0(n1423), .B0(n1240), .CO(n1238), .S0(n1267) );
  HS65_GSS_XOR3X2 U1331 ( .A(x_z2[5]), .B(n1268), .C(n1267), .Z(
        \mul_b1/fa1_s1[15] ) );
  HS65_GS_HA1X4 U1332 ( .A0(n1421), .B0(n1241), .CO(n1240), .S0(n1270) );
  HS65_GS_HA1X4 U1333 ( .A0(n1425), .B0(n1242), .CO(n1239), .S0(n1269) );
  HS65_GSS_XOR3X2 U1334 ( .A(x_z2[4]), .B(n1270), .C(n1269), .Z(
        \mul_b1/fa1_s1[14] ) );
  HS65_GS_HA1X4 U1335 ( .A0(n1423), .B0(n1243), .CO(n1242), .S0(n1272) );
  HS65_GS_HA1X4 U1336 ( .A0(n1419), .B0(n1244), .CO(n1241), .S0(n1271) );
  HS65_GSS_XOR3X2 U1337 ( .A(x_z2[3]), .B(n1272), .C(n1271), .Z(
        \mul_b1/fa1_s1[13] ) );
  HS65_GS_HA1X4 U1338 ( .A0(n1418), .B0(n1245), .CO(n1244), .S0(n1274) );
  HS65_GS_HA1X4 U1339 ( .A0(n1421), .B0(n1246), .CO(n1243), .S0(n1273) );
  HS65_GSS_XOR3X2 U1340 ( .A(x_z2[2]), .B(n1274), .C(n1273), .Z(
        \mul_b1/fa1_s1[12] ) );
  HS65_GS_HA1X4 U1341 ( .A0(n1419), .B0(n1247), .CO(n1246), .S0(n1276) );
  HS65_GS_HA1X4 U1342 ( .A0(n1416), .B0(n1248), .CO(n1245), .S0(n1275) );
  HS65_GSS_XOR3X2 U1343 ( .A(x_z2[1]), .B(n1276), .C(n1275), .Z(
        \mul_b1/fa1_s1[11] ) );
  HS65_GS_HA1X4 U1344 ( .A0(n1418), .B0(n1249), .CO(n1247), .S0(n1278) );
  HS65_GS_HA1X4 U1345 ( .A0(n1414), .B0(n1250), .CO(n1248), .S0(n1277) );
  HS65_GSS_XOR3X2 U1346 ( .A(x_z2[0]), .B(n1278), .C(n1277), .Z(
        \mul_b1/fa1_s1[10] ) );
  HS65_GS_HA1X4 U1347 ( .A0(n1416), .B0(n1251), .CO(n1249), .S0(n1280) );
  HS65_GS_HA1X4 U1348 ( .A0(n1752), .B0(n1411), .CO(n1250), .S0(n1279) );
  HS65_GSS_XOR2X3 U1349 ( .A(n1280), .B(n1279), .Z(\mul_b1/fa1_s1[9] ) );
  HS65_GS_HA1X4 U1350 ( .A0(n1414), .B0(n1252), .CO(n1251), .S0(n1281) );
  HS65_GSS_XOR2X3 U1351 ( .A(n1281), .B(x_z2[0]), .Z(\mul_b1/fa1_s1[8] ) );
  HS65_GS_PAO2X4 U1352 ( .A(n1254), .B(n1253), .P(x_z2[12]), .Z(
        \mul_b1/fa1_c1[22] ) );
  HS65_GS_PAO2X4 U1353 ( .A(n1256), .B(n1255), .P(x_z2[11]), .Z(
        \mul_b1/fa1_c1[21] ) );
  HS65_GS_PAO2X4 U1354 ( .A(n1258), .B(n1257), .P(x_z2[10]), .Z(
        \mul_b1/fa1_c1[20] ) );
  HS65_GS_PAO2X4 U1355 ( .A(n1260), .B(n1259), .P(x_z2[9]), .Z(
        \mul_b1/fa1_c1[19] ) );
  HS65_GS_PAO2X4 U1356 ( .A(n1262), .B(n1261), .P(x_z2[8]), .Z(
        \mul_b1/fa1_c1[18] ) );
  HS65_GS_PAO2X4 U1357 ( .A(n1264), .B(n1263), .P(x_z2[7]), .Z(
        \mul_b1/fa1_c1[17] ) );
  HS65_GS_PAO2X4 U1358 ( .A(n1266), .B(n1265), .P(x_z2[6]), .Z(
        \mul_b1/fa1_c1[16] ) );
  HS65_GS_PAO2X4 U1359 ( .A(n1268), .B(n1267), .P(x_z2[5]), .Z(
        \mul_b1/fa1_c1[15] ) );
  HS65_GS_PAO2X4 U1360 ( .A(n1270), .B(n1269), .P(x_z2[4]), .Z(
        \mul_b1/fa1_c1[14] ) );
  HS65_GS_PAO2X4 U1361 ( .A(n1272), .B(n1271), .P(x_z2[3]), .Z(
        \mul_b1/fa1_c1[13] ) );
  HS65_GS_PAO2X4 U1362 ( .A(n1274), .B(n1273), .P(x_z2[2]), .Z(
        \mul_b1/fa1_c1[12] ) );
  HS65_GS_PAO2X4 U1363 ( .A(n1276), .B(n1275), .P(x_z2[1]), .Z(
        \mul_b1/fa1_c1[11] ) );
  HS65_GS_PAO2X4 U1364 ( .A(n1278), .B(n1277), .P(x_z2[0]), .Z(
        \mul_b1/fa1_c1[10] ) );
  HS65_GS_AND2X4 U1365 ( .A(n1280), .B(n1279), .Z(\mul_b1/fa1_c1[9] ) );
  HS65_GS_AND2X4 U1366 ( .A(n1281), .B(x_z2[0]), .Z(\mul_b1/fa1_c1[8] ) );
  HS65_GS_NOR2X2 U1367 ( .A(\DP_OP_331J1_157_5454/n87 ), .B(n1282), .Z(n1283)
         );
  HS65_GSS_XNOR2X3 U1368 ( .A(n1283), .B(n1439), .Z(\mul_b1/fa1_s2[29] ) );
  HS65_GS_HA1X4 U1369 ( .A0(n1700), .B0(n1284), .CO(n1296), .S0(n1310) );
  HS65_GSS_XNOR2X3 U1370 ( .A(y_z2[15]), .B(n1441), .Z(n1297) );
  HS65_GSS_XNOR2X3 U1371 ( .A(n1297), .B(n1676), .Z(\mul_a2/fa1_s0[16] ) );
  HS65_GS_HA1X4 U1372 ( .A0(n1676), .B0(n1285), .CO(n1441), .S0(n1298) );
  HS65_GSS_XNOR2X3 U1373 ( .A(n1298), .B(n1678), .Z(\mul_a2/fa1_s0[15] ) );
  HS65_GS_HA1X4 U1374 ( .A0(n1678), .B0(n1286), .CO(n1285), .S0(n1299) );
  HS65_GSS_XNOR2X3 U1375 ( .A(n1299), .B(n1680), .Z(\mul_a2/fa1_s0[14] ) );
  HS65_GS_HA1X4 U1376 ( .A0(n1680), .B0(n1287), .CO(n1286), .S0(n1300) );
  HS65_GSS_XNOR2X3 U1377 ( .A(n1300), .B(n1682), .Z(\mul_a2/fa1_s0[13] ) );
  HS65_GS_HA1X4 U1378 ( .A0(n1682), .B0(n1288), .CO(n1287), .S0(n1301) );
  HS65_GSS_XNOR2X3 U1379 ( .A(n1301), .B(n1684), .Z(\mul_a2/fa1_s0[12] ) );
  HS65_GS_HA1X4 U1380 ( .A0(n1684), .B0(n1289), .CO(n1288), .S0(n1302) );
  HS65_GSS_XNOR2X3 U1381 ( .A(n1302), .B(n1686), .Z(\mul_a2/fa1_s0[11] ) );
  HS65_GS_HA1X4 U1382 ( .A0(n1686), .B0(n1290), .CO(n1289), .S0(n1303) );
  HS65_GSS_XNOR2X3 U1383 ( .A(n1303), .B(n1688), .Z(\mul_a2/fa1_s0[10] ) );
  HS65_GS_HA1X4 U1384 ( .A0(n1688), .B0(n1291), .CO(n1290), .S0(n1304) );
  HS65_GSS_XNOR2X3 U1385 ( .A(n1304), .B(n1690), .Z(\mul_a2/fa1_s0[9] ) );
  HS65_GS_HA1X4 U1386 ( .A0(n1690), .B0(n1292), .CO(n1291), .S0(n1305) );
  HS65_GSS_XNOR2X3 U1387 ( .A(n1305), .B(n1692), .Z(\mul_a2/fa1_s0[8] ) );
  HS65_GS_HA1X4 U1388 ( .A0(n1692), .B0(n1293), .CO(n1292), .S0(n1306) );
  HS65_GSS_XNOR2X3 U1389 ( .A(n1306), .B(n1694), .Z(\mul_a2/fa1_s0[7] ) );
  HS65_GS_HA1X4 U1390 ( .A0(n1694), .B0(n1294), .CO(n1293), .S0(n1307) );
  HS65_GSS_XNOR2X3 U1391 ( .A(n1307), .B(n1696), .Z(\mul_a2/fa1_s0[6] ) );
  HS65_GS_HA1X4 U1392 ( .A0(n1696), .B0(n1295), .CO(n1294), .S0(n1308) );
  HS65_GSS_XNOR2X3 U1393 ( .A(n1308), .B(n1698), .Z(\mul_a2/fa1_s0[5] ) );
  HS65_GS_HA1X4 U1394 ( .A0(n1698), .B0(n1296), .CO(n1295), .S0(n1309) );
  HS65_GSS_XNOR2X3 U1395 ( .A(n1309), .B(n1700), .Z(\mul_a2/fa1_s0[4] ) );
  HS65_GS_AND2X4 U1396 ( .A(y_z2[14]), .B(n1297), .Z(\mul_a2/fa1_c0[16] ) );
  HS65_GS_AND2X4 U1397 ( .A(n1298), .B(y_z2[13]), .Z(\mul_a2/fa1_c0[15] ) );
  HS65_GS_AND2X4 U1398 ( .A(y_z2[12]), .B(n1299), .Z(\mul_a2/fa1_c0[14] ) );
  HS65_GS_AND2X4 U1399 ( .A(y_z2[11]), .B(n1300), .Z(\mul_a2/fa1_c0[13] ) );
  HS65_GS_AND2X4 U1400 ( .A(n1301), .B(y_z2[10]), .Z(\mul_a2/fa1_c0[12] ) );
  HS65_GS_AND2X4 U1401 ( .A(n1302), .B(y_z2[9]), .Z(\mul_a2/fa1_c0[11] ) );
  HS65_GS_AND2X4 U1402 ( .A(y_z2[8]), .B(n1303), .Z(\mul_a2/fa1_c0[10] ) );
  HS65_GS_AND2X4 U1403 ( .A(y_z2[7]), .B(n1304), .Z(\mul_a2/fa1_c0[9] ) );
  HS65_GS_AND2X4 U1404 ( .A(y_z2[6]), .B(n1305), .Z(\mul_a2/fa1_c0[8] ) );
  HS65_GS_AND2X4 U1405 ( .A(y_z2[5]), .B(n1306), .Z(\mul_a2/fa1_c0[7] ) );
  HS65_GS_AND2X4 U1406 ( .A(y_z2[4]), .B(n1307), .Z(\mul_a2/fa1_c0[6] ) );
  HS65_GS_AND2X4 U1407 ( .A(y_z2[3]), .B(n1308), .Z(\mul_a2/fa1_c0[5] ) );
  HS65_GS_AND2X4 U1408 ( .A(y_z2[2]), .B(n1309), .Z(\mul_a2/fa1_c0[4] ) );
  HS65_GS_AND2X4 U1409 ( .A(n1310), .B(y_z2[1]), .Z(\mul_a2/fa1_c0[3] ) );
  HS65_GS_HA1X4 U1410 ( .A0(n1702), .B0(n1701), .CO(n1284), .S0(n1311) );
  HS65_GS_AND2X4 U1411 ( .A(n1311), .B(y_z2[0]), .Z(\mul_a2/fa1_c0[2] ) );
  HS65_GS_FA1X4 U1412 ( .A0(n1314), .B0(n1313), .CI(n1312), .CO(n672), .S0(
        n1315) );
  HS65_GS_AO12X4 U1413 ( .A(n1315), .B(n1341), .C(n1340), .Z(
        \mul_a2/result_sat[12] ) );
  HS65_GS_FA1X4 U1414 ( .A0(n1318), .B0(n1317), .CI(n1316), .CO(n1314), .S0(
        n1319) );
  HS65_GS_AO12X4 U1415 ( .A(n1319), .B(n1341), .C(n1340), .Z(
        \mul_a2/result_sat[11] ) );
  HS65_GS_FA1X4 U1416 ( .A0(n1322), .B0(n1321), .CI(n1320), .CO(n1318), .S0(
        n1323) );
  HS65_GS_AO12X4 U1417 ( .A(n1323), .B(n1341), .C(n1340), .Z(
        \mul_a2/result_sat[10] ) );
  HS65_GS_FA1X4 U1418 ( .A0(n1326), .B0(n1325), .CI(n1324), .CO(n1322), .S0(
        n1327) );
  HS65_GS_AO12X4 U1419 ( .A(n1327), .B(n1341), .C(n1340), .Z(
        \mul_a2/result_sat[9] ) );
  HS65_GS_FA1X4 U1420 ( .A0(n1330), .B0(n1329), .CI(n1328), .CO(n1324), .S0(
        n1331) );
  HS65_GS_OA12X4 U1421 ( .A(n1340), .B(n1331), .C(n1341), .Z(
        \mul_a2/result_sat[8] ) );
  HS65_GS_FA1X4 U1422 ( .A0(n1334), .B0(n1333), .CI(n1332), .CO(n1328), .S0(
        n1335) );
  HS65_GS_AO12X4 U1423 ( .A(n1335), .B(n1341), .C(n1340), .Z(
        \mul_a2/result_sat[7] ) );
  HS65_GS_FA1X4 U1424 ( .A0(n1338), .B0(n1337), .CI(n1336), .CO(n1332), .S0(
        n1339) );
  HS65_GS_OA12X4 U1425 ( .A(n1340), .B(n1339), .C(n1341), .Z(
        \mul_a2/result_sat[6] ) );
  HS65_GS_IVX2 U1426 ( .A(n1341), .Z(n1762) );
  HS65_GS_OAI21X2 U1427 ( .A(n1344), .B(n1343), .C(n1342), .Z(n1345) );
  HS65_GS_OAI21X2 U1428 ( .A(n1762), .B(n1345), .C(n1763), .Z(
        \mul_a2/result_sat[3] ) );
  HS65_GS_OAI21X2 U1429 ( .A(n1347), .B(n1346), .C(n1757), .Z(n1348) );
  HS65_GS_OAI21X2 U1430 ( .A(n1762), .B(n1348), .C(n1763), .Z(
        \mul_a2/result_sat[0] ) );
  HS65_GS_MUX21X4 U1431 ( .D0(y_z1[1]), .D1(data_out[1]), .S0(n1821), .Z(n1913) );
  HS65_GS_IVX2 U1432 ( .A(n1448), .Z(n1404) );
  HS65_GS_OAI112X1 U1433 ( .A(n1350), .B(p_a1[1]), .C(n1403), .D(n1349), .Z(
        n1351) );
  HS65_GS_AO22X4 U1434 ( .A(data_out[1]), .B(n1810), .C(n1404), .D(n1351), .Z(
        n1912) );
  HS65_GS_MUXI21X2 U1435 ( .D0(n1700), .D1(n1754), .S0(n1437), .Z(n1911) );
  HS65_GS_OAI112X1 U1436 ( .A(n1354), .B(n1353), .C(n1403), .D(n1352), .Z(
        n1355) );
  HS65_GS_AO22X4 U1437 ( .A(data_out[2]), .B(n1810), .C(n1404), .D(n1355), .Z(
        n1909) );
  HS65_GS_MUXI21X2 U1438 ( .D0(n1698), .D1(n1720), .S0(n1437), .Z(n1908) );
  HS65_GS_AOI112X2 U1439 ( .A(n1358), .B(n1357), .C(n1448), .D(n1356), .Z(
        n1359) );
  HS65_GS_IVX2 U1440 ( .A(n1403), .Z(n1445) );
  HS65_GS_AO112X4 U1441 ( .A(data_out[3]), .B(n1810), .C(n1359), .D(n1445), 
        .Z(n1906) );
  HS65_GS_MUXI21X2 U1442 ( .D0(n1696), .D1(n1718), .S0(n1437), .Z(n1905) );
  HS65_GS_IVX2 U1443 ( .A(data_out[4]), .Z(n1366) );
  HS65_GS_MUXI21X2 U1444 ( .D0(n1718), .D1(n1366), .S0(valid_in), .Z(n1904) );
  HS65_GSS_XOR2X3 U1445 ( .A(n1361), .B(n1360), .Z(n1364) );
  HS65_GS_OAI21X2 U1446 ( .A(n1363), .B(n1364), .C(n1403), .Z(n1362) );
  HS65_GS_CBI4I1X3 U1447 ( .A(n1364), .B(n1363), .C(n1362), .D(n1404), .Z(
        n1365) );
  HS65_GS_OAI21X2 U1448 ( .A(valid_T3), .B(n1366), .C(n1365), .Z(n1903) );
  HS65_GS_MUXI21X2 U1449 ( .D0(n1694), .D1(n1716), .S0(n1437), .Z(n1902) );
  HS65_GS_IVX2 U1450 ( .A(data_out[5]), .Z(n1371) );
  HS65_GS_MUXI21X2 U1451 ( .D0(n1716), .D1(n1371), .S0(valid_in), .Z(n1901) );
  HS65_GS_OAI21X2 U1452 ( .A(n1368), .B(n1369), .C(n1403), .Z(n1367) );
  HS65_GS_CBI4I1X3 U1453 ( .A(n1369), .B(n1368), .C(n1367), .D(n1404), .Z(
        n1370) );
  HS65_GS_OAI21X2 U1454 ( .A(valid_T3), .B(n1371), .C(n1370), .Z(n1900) );
  HS65_GS_MUXI21X2 U1455 ( .D0(n1692), .D1(n1740), .S0(valid_in), .Z(n1899) );
  HS65_GS_FA1X4 U1456 ( .A0(n1374), .B0(n1373), .CI(n1372), .CO(n766), .S0(
        n1376) );
  HS65_GS_AOI12X2 U1457 ( .A(data_out[6]), .B(n1810), .C(n1445), .Z(n1375) );
  HS65_GS_OAI21X2 U1458 ( .A(n1448), .B(n1376), .C(n1375), .Z(n1897) );
  HS65_GS_MUXI21X2 U1459 ( .D0(n1690), .D1(n1738), .S0(n1821), .Z(n1896) );
  HS65_GS_MUXI21X2 U1460 ( .D0(n1688), .D1(n1736), .S0(n1821), .Z(n1893) );
  HS65_GS_MUXI21X2 U1461 ( .D0(n1686), .D1(n1734), .S0(valid_in), .Z(n1890) );
  HS65_GS_IVX2 U1462 ( .A(data_out[9]), .Z(n1383) );
  HS65_GS_MUXI21X2 U1463 ( .D0(n1734), .D1(n1383), .S0(n1821), .Z(n1889) );
  HS65_GSS_XOR2X3 U1464 ( .A(n1378), .B(n1377), .Z(n1381) );
  HS65_GS_OAI21X2 U1465 ( .A(n1380), .B(n1381), .C(n1403), .Z(n1379) );
  HS65_GS_CBI4I1X3 U1466 ( .A(n1381), .B(n1380), .C(n1379), .D(n1404), .Z(
        n1382) );
  HS65_GS_OAI21X2 U1467 ( .A(valid_T3), .B(n1383), .C(n1382), .Z(n1888) );
  HS65_GS_MUXI21X2 U1468 ( .D0(n1684), .D1(n1732), .S0(n1821), .Z(n1887) );
  HS65_GS_OAI112X1 U1469 ( .A(n1386), .B(n1385), .C(n1403), .D(n1384), .Z(
        n1387) );
  HS65_GS_AO22X4 U1470 ( .A(data_out[10]), .B(n1810), .C(n1404), .D(n1387), 
        .Z(n1885) );
  HS65_GS_MUXI21X2 U1471 ( .D0(n1682), .D1(n1730), .S0(valid_in), .Z(n1884) );
  HS65_GS_OAI112X1 U1472 ( .A(n1390), .B(n1389), .C(n1403), .D(n1388), .Z(
        n1391) );
  HS65_GS_AO22X4 U1473 ( .A(data_out[11]), .B(n1810), .C(n1404), .D(n1391), 
        .Z(n1882) );
  HS65_GS_MUXI21X2 U1474 ( .D0(n1680), .D1(n1728), .S0(n1821), .Z(n1881) );
  HS65_GS_OAI112X1 U1475 ( .A(n1394), .B(n1393), .C(n1403), .D(n1392), .Z(
        n1395) );
  HS65_GS_AO22X4 U1476 ( .A(data_out[12]), .B(n1810), .C(n1404), .D(n1395), 
        .Z(n1879) );
  HS65_GS_MUXI21X2 U1477 ( .D0(n1678), .D1(n1726), .S0(valid_in), .Z(n1878) );
  HS65_GS_IVX2 U1478 ( .A(data_out[13]), .Z(n1402) );
  HS65_GS_MUXI21X2 U1479 ( .D0(n1726), .D1(n1402), .S0(valid_in), .Z(n1877) );
  HS65_GSS_XOR2X3 U1480 ( .A(n1397), .B(n1396), .Z(n1400) );
  HS65_GS_OAI21X2 U1481 ( .A(n1399), .B(n1400), .C(n1403), .Z(n1398) );
  HS65_GS_CBI4I1X3 U1482 ( .A(n1400), .B(n1399), .C(n1398), .D(n1404), .Z(
        n1401) );
  HS65_GS_OAI21X2 U1483 ( .A(valid_T3), .B(n1402), .C(n1401), .Z(n1876) );
  HS65_GS_MUXI21X2 U1484 ( .D0(n1676), .D1(n1724), .S0(n1821), .Z(n1875) );
  HS65_GS_IVX2 U1485 ( .A(data_out[14]), .Z(n1409) );
  HS65_GS_MUXI21X2 U1486 ( .D0(n1724), .D1(n1409), .S0(valid_in), .Z(n1874) );
  HS65_GS_OAI21X2 U1487 ( .A(n1406), .B(n1407), .C(n1403), .Z(n1405) );
  HS65_GS_CBI4I1X3 U1488 ( .A(n1407), .B(n1406), .C(n1405), .D(n1404), .Z(
        n1408) );
  HS65_GS_OAI21X2 U1489 ( .A(valid_T3), .B(n1409), .C(n1408), .Z(n1873) );
  HS65_GS_IVX2 U1490 ( .A(y_z2[15]), .Z(n1442) );
  HS65_GS_MUXI21X2 U1491 ( .D0(n1442), .D1(n1705), .S0(valid_in), .Z(n1872) );
  HS65_GS_IVX2 U1492 ( .A(data_out[15]), .Z(n1809) );
  HS65_GS_MUXI21X2 U1493 ( .D0(n1705), .D1(n1809), .S0(n1821), .Z(n1871) );
  HS65_GS_MUXI21X2 U1494 ( .D0(n1741), .D1(n1411), .S0(valid_in), .Z(n1869) );
  HS65_GS_MUXI21X2 U1495 ( .D0(n1411), .D1(n1410), .S0(n1821), .Z(n1868) );
  HS65_GS_MUXI21X2 U1496 ( .D0(n1742), .D1(n1752), .S0(n1437), .Z(n1867) );
  HS65_GS_BFX4 U1497 ( .A(valid_in), .Z(n1434) );
  HS65_GS_MUXI21X2 U1498 ( .D0(n1752), .D1(n1412), .S0(n1434), .Z(n1866) );
  HS65_GS_MUXI21X2 U1499 ( .D0(n1751), .D1(n1414), .S0(valid_in), .Z(n1865) );
  HS65_GS_MUXI21X2 U1500 ( .D0(n1414), .D1(n1413), .S0(n1821), .Z(n1864) );
  HS65_GS_MUXI21X2 U1501 ( .D0(n1518), .D1(n1416), .S0(n1437), .Z(n1863) );
  HS65_GS_MUXI21X2 U1502 ( .D0(n1416), .D1(n1415), .S0(n1434), .Z(n1862) );
  HS65_GS_MUXI21X2 U1503 ( .D0(n1516), .D1(n1418), .S0(valid_in), .Z(n1861) );
  HS65_GS_MUXI21X2 U1504 ( .D0(n1418), .D1(n1417), .S0(n1440), .Z(n1860) );
  HS65_GS_MUX21X4 U1505 ( .D0(y_z2[1]), .D1(y_z1[1]), .S0(n1821), .Z(n1914) );
  HS65_GS_MUXI21X2 U1506 ( .D0(n1514), .D1(n1419), .S0(n1437), .Z(n1859) );
  HS65_GS_MUXI21X2 U1507 ( .D0(n1419), .D1(n1420), .S0(n1437), .Z(n1858) );
  HS65_GS_MUXI21X2 U1508 ( .D0(n1512), .D1(n1421), .S0(n1437), .Z(n1857) );
  HS65_GS_MUXI21X2 U1509 ( .D0(n1421), .D1(n1422), .S0(n1437), .Z(n1856) );
  HS65_GS_MUXI21X2 U1510 ( .D0(n1510), .D1(n1423), .S0(n1434), .Z(n1855) );
  HS65_GS_MUXI21X2 U1511 ( .D0(n1423), .D1(n1424), .S0(n1434), .Z(n1854) );
  HS65_GS_MUXI21X2 U1512 ( .D0(n1508), .D1(n1425), .S0(n1434), .Z(n1853) );
  HS65_GS_MUXI21X2 U1513 ( .D0(n1425), .D1(n1426), .S0(n1434), .Z(n1852) );
  HS65_GS_MUXI21X2 U1514 ( .D0(n1506), .D1(n1428), .S0(n1440), .Z(n1851) );
  HS65_GS_MUXI21X2 U1515 ( .D0(n1428), .D1(n1427), .S0(n1434), .Z(n1850) );
  HS65_GS_MUXI21X2 U1516 ( .D0(n1504), .D1(n1429), .S0(n1434), .Z(n1849) );
  HS65_GS_MUXI21X2 U1517 ( .D0(n1429), .D1(n1430), .S0(n1434), .Z(n1848) );
  HS65_GS_MUXI21X2 U1518 ( .D0(n1502), .D1(n1432), .S0(n1434), .Z(n1847) );
  HS65_GS_MUXI21X2 U1519 ( .D0(n1432), .D1(n1431), .S0(n1434), .Z(n1846) );
  HS65_GS_MUXI21X2 U1520 ( .D0(n1500), .D1(n1749), .S0(n1434), .Z(n1845) );
  HS65_GS_MUXI21X2 U1521 ( .D0(n1749), .D1(n1433), .S0(n1434), .Z(n1844) );
  HS65_GS_MUXI21X2 U1522 ( .D0(n1498), .D1(n1747), .S0(n1434), .Z(n1843) );
  HS65_GS_MUXI21X2 U1523 ( .D0(n1747), .D1(n1435), .S0(n1434), .Z(n1842) );
  HS65_GS_MUXI21X2 U1524 ( .D0(n1496), .D1(n1745), .S0(n1437), .Z(n1841) );
  HS65_GS_MUXI21X2 U1525 ( .D0(n1745), .D1(n1436), .S0(n1437), .Z(n1840) );
  HS65_GS_MUXI21X2 U1526 ( .D0(n1494), .D1(n1439), .S0(n1437), .Z(n1839) );
  HS65_GS_MUXI21X2 U1527 ( .D0(n1439), .D1(n1438), .S0(n1437), .Z(n1838) );
  HS65_GS_MUX21X4 U1528 ( .D0(x_z1[0]), .D1(data_in[0]), .S0(n1821), .Z(n1837)
         );
  HS65_GS_MUX21X4 U1529 ( .D0(x_z1[1]), .D1(data_in[1]), .S0(n1821), .Z(n1836)
         );
  HS65_GS_MUX21X4 U1530 ( .D0(x_z1[2]), .D1(data_in[2]), .S0(n1821), .Z(n1835)
         );
  HS65_GS_MUX21X4 U1531 ( .D0(x_z1[3]), .D1(data_in[3]), .S0(n1821), .Z(n1834)
         );
  HS65_GS_MUX21X4 U1532 ( .D0(x_z1[4]), .D1(data_in[4]), .S0(n1821), .Z(n1833)
         );
  HS65_GS_MUX21X4 U1533 ( .D0(x_z1[5]), .D1(data_in[5]), .S0(n1440), .Z(n1832)
         );
  HS65_GS_MUX21X4 U1534 ( .D0(x_z1[6]), .D1(data_in[6]), .S0(n1440), .Z(n1831)
         );
  HS65_GS_MUX21X4 U1535 ( .D0(x_z1[7]), .D1(data_in[7]), .S0(n1440), .Z(n1830)
         );
  HS65_GS_MUX21X4 U1536 ( .D0(x_z1[8]), .D1(data_in[8]), .S0(n1440), .Z(n1829)
         );
  HS65_GS_MUX21X4 U1537 ( .D0(x_z1[9]), .D1(data_in[9]), .S0(n1440), .Z(n1828)
         );
  HS65_GS_MUX21X4 U1538 ( .D0(x_z1[10]), .D1(data_in[10]), .S0(n1440), .Z(
        n1827) );
  HS65_GS_MUX21X4 U1539 ( .D0(x_z1[11]), .D1(data_in[11]), .S0(n1440), .Z(
        n1826) );
  HS65_GS_MUX21X4 U1540 ( .D0(x_z1[12]), .D1(data_in[12]), .S0(n1821), .Z(
        n1825) );
  HS65_GS_MUX21X4 U1541 ( .D0(x_z1[13]), .D1(data_in[13]), .S0(n1440), .Z(
        n1824) );
  HS65_GS_MUX21X4 U1542 ( .D0(x_z1[14]), .D1(data_in[14]), .S0(n1440), .Z(
        n1823) );
  HS65_GS_MUX21X4 U1543 ( .D0(n1820), .D1(data_in[15]), .S0(n1821), .Z(n1822)
         );
  HS65_GS_NOR2X2 U1544 ( .A(y_z2[15]), .B(n1441), .Z(n1443) );
  HS65_GSS_XNOR2X6 U1545 ( .A(n1443), .B(n1442), .Z(\mul_a2/fa1_s0[31] ) );
  HS65_GS_FA1X4 U1546 ( .A0(p_a2[0]), .B0(p_a1[0]), .CI(n1444), .CO(n712), 
        .S0(n1447) );
  HS65_GS_AOI12X2 U1547 ( .A(data_out[0]), .B(n1810), .C(n1445), .Z(n1446) );
  HS65_GS_OAI21X2 U1548 ( .A(n1448), .B(n1447), .C(n1446), .Z(n1915) );
  HS65_GSS_XNOR2X3 U1549 ( .A(\DP_OP_371J1_181_1383/n79 ), .B(n1449), .Z(n1659) );
  HS65_GS_IVX2 U1550 ( .A(n1659), .Z(n1450) );
  HS65_GS_OAI21X2 U1551 ( .A(n1494), .B(n1450), .C(n1496), .Z(
        \mul_b2/fa1_c0[18] ) );
  HS65_GS_HA1X4 U1552 ( .A0(n1496), .B0(n1451), .CO(n1449), .S0(n1660) );
  HS65_GS_IVX2 U1553 ( .A(n1660), .Z(n1453) );
  HS65_GS_OAI21X2 U1554 ( .A(\DP_OP_371J1_181_1383/n79 ), .B(n1660), .C(
        x_reg2[13]), .Z(n1452) );
  HS65_GS_OAI21X2 U1555 ( .A(n1494), .B(n1453), .C(n1452), .Z(
        \mul_b2/fa1_c0[17] ) );
  HS65_GS_HA1X4 U1556 ( .A0(n1498), .B0(n1454), .CO(n1451), .S0(n1661) );
  HS65_GS_IVX2 U1557 ( .A(n1661), .Z(n1456) );
  HS65_GS_OAI21X2 U1558 ( .A(\DP_OP_371J1_181_1383/n79 ), .B(n1661), .C(
        x_reg2[12]), .Z(n1455) );
  HS65_GS_OAI21X2 U1559 ( .A(n1494), .B(n1456), .C(n1455), .Z(
        \mul_b2/fa1_c0[16] ) );
  HS65_GS_HA1X4 U1560 ( .A0(n1500), .B0(n1457), .CO(n1454), .S0(n1662) );
  HS65_GS_IVX2 U1561 ( .A(n1662), .Z(n1459) );
  HS65_GS_OAI21X2 U1562 ( .A(\DP_OP_371J1_181_1383/n79 ), .B(n1662), .C(
        x_reg2[11]), .Z(n1458) );
  HS65_GS_OAI21X2 U1563 ( .A(n1494), .B(n1459), .C(n1458), .Z(
        \mul_b2/fa1_c0[15] ) );
  HS65_GS_HA1X4 U1564 ( .A0(n1502), .B0(n1460), .CO(n1457), .S0(n1663) );
  HS65_GS_IVX2 U1565 ( .A(n1663), .Z(n1462) );
  HS65_GS_OAI21X2 U1566 ( .A(x_reg2[14]), .B(n1663), .C(x_reg2[10]), .Z(n1461)
         );
  HS65_GS_OAI21X2 U1567 ( .A(n1496), .B(n1462), .C(n1461), .Z(
        \mul_b2/fa1_c0[14] ) );
  HS65_GS_HA1X4 U1568 ( .A0(n1504), .B0(n1463), .CO(n1460), .S0(n1664) );
  HS65_GS_IVX2 U1569 ( .A(n1664), .Z(n1465) );
  HS65_GS_OAI21X2 U1570 ( .A(x_reg2[13]), .B(n1664), .C(x_reg2[9]), .Z(n1464)
         );
  HS65_GS_OAI21X2 U1571 ( .A(n1498), .B(n1465), .C(n1464), .Z(
        \mul_b2/fa1_c0[13] ) );
  HS65_GS_HA1X4 U1572 ( .A0(n1506), .B0(n1466), .CO(n1463), .S0(n1665) );
  HS65_GS_IVX2 U1573 ( .A(n1665), .Z(n1468) );
  HS65_GS_OAI21X2 U1574 ( .A(x_reg2[12]), .B(n1665), .C(x_reg2[8]), .Z(n1467)
         );
  HS65_GS_OAI21X2 U1575 ( .A(n1500), .B(n1468), .C(n1467), .Z(
        \mul_b2/fa1_c0[12] ) );
  HS65_GS_HA1X4 U1576 ( .A0(n1508), .B0(n1469), .CO(n1466), .S0(n1666) );
  HS65_GS_IVX2 U1577 ( .A(n1666), .Z(n1471) );
  HS65_GS_OAI21X2 U1578 ( .A(x_reg2[11]), .B(n1666), .C(x_reg2[7]), .Z(n1470)
         );
  HS65_GS_OAI21X2 U1579 ( .A(n1502), .B(n1471), .C(n1470), .Z(
        \mul_b2/fa1_c0[11] ) );
  HS65_GS_HA1X4 U1580 ( .A0(n1510), .B0(n1472), .CO(n1469), .S0(n1667) );
  HS65_GS_IVX2 U1581 ( .A(n1667), .Z(n1474) );
  HS65_GS_OAI21X2 U1582 ( .A(x_reg2[10]), .B(n1667), .C(x_reg2[6]), .Z(n1473)
         );
  HS65_GS_OAI21X2 U1583 ( .A(n1504), .B(n1474), .C(n1473), .Z(
        \mul_b2/fa1_c0[10] ) );
  HS65_GS_HA1X4 U1584 ( .A0(n1512), .B0(n1475), .CO(n1472), .S0(n1668) );
  HS65_GS_IVX2 U1585 ( .A(n1668), .Z(n1477) );
  HS65_GS_OAI21X2 U1586 ( .A(x_reg2[9]), .B(n1668), .C(x_reg2[5]), .Z(n1476)
         );
  HS65_GS_OAI21X2 U1587 ( .A(n1506), .B(n1477), .C(n1476), .Z(
        \mul_b2/fa1_c0[9] ) );
  HS65_GS_HA1X4 U1588 ( .A0(n1514), .B0(n1478), .CO(n1475), .S0(n1669) );
  HS65_GS_IVX2 U1589 ( .A(n1669), .Z(n1480) );
  HS65_GS_OAI21X2 U1590 ( .A(x_reg2[8]), .B(n1669), .C(x_reg2[4]), .Z(n1479)
         );
  HS65_GS_OAI21X2 U1591 ( .A(n1508), .B(n1480), .C(n1479), .Z(
        \mul_b2/fa1_c0[8] ) );
  HS65_GS_HA1X4 U1592 ( .A0(n1516), .B0(n1481), .CO(n1478), .S0(n1670) );
  HS65_GS_IVX2 U1593 ( .A(n1670), .Z(n1483) );
  HS65_GS_OAI21X2 U1594 ( .A(x_reg2[7]), .B(n1670), .C(x_reg2[3]), .Z(n1482)
         );
  HS65_GS_OAI21X2 U1595 ( .A(n1510), .B(n1483), .C(n1482), .Z(
        \mul_b2/fa1_c0[7] ) );
  HS65_GS_HA1X4 U1596 ( .A0(n1518), .B0(n1484), .CO(n1481), .S0(n1671) );
  HS65_GS_IVX2 U1597 ( .A(n1671), .Z(n1486) );
  HS65_GS_OAI21X2 U1598 ( .A(x_reg2[6]), .B(n1671), .C(x_reg2[2]), .Z(n1485)
         );
  HS65_GS_OAI21X2 U1599 ( .A(n1512), .B(n1486), .C(n1485), .Z(
        \mul_b2/fa1_c0[6] ) );
  HS65_GS_HA1X4 U1600 ( .A0(n1751), .B0(n1487), .CO(n1484), .S0(n1672) );
  HS65_GS_IVX2 U1601 ( .A(n1672), .Z(n1489) );
  HS65_GS_OAI21X2 U1602 ( .A(x_reg2[5]), .B(n1672), .C(x_reg2[1]), .Z(n1488)
         );
  HS65_GS_OAI21X2 U1603 ( .A(n1514), .B(n1489), .C(n1488), .Z(
        \mul_b2/fa1_c0[5] ) );
  HS65_GS_HA1X4 U1604 ( .A0(n1742), .B0(n1741), .CO(n1487), .S0(n1673) );
  HS65_GS_IVX2 U1605 ( .A(n1673), .Z(n1491) );
  HS65_GS_OAI21X2 U1606 ( .A(x_reg2[4]), .B(n1673), .C(x_reg2[0]), .Z(n1490)
         );
  HS65_GS_OAI21X2 U1607 ( .A(n1516), .B(n1491), .C(n1490), .Z(
        \mul_b2/fa1_c0[4] ) );
  HS65_GS_AND2X4 U1608 ( .A(x_reg2[3]), .B(x_reg2[0]), .Z(\mul_b2/fa1_c0[3] )
         );
  HS65_GSS_XNOR2X3 U1609 ( .A(n1519), .B(n1496), .Z(\mul_b2/fa1_s1[23] ) );
  HS65_GSS_XNOR2X3 U1610 ( .A(\DP_OP_371J1_181_1383/n79 ), .B(n1492), .Z(n1520) );
  HS65_GSS_XNOR2X3 U1611 ( .A(n1520), .B(n1498), .Z(\mul_b2/fa1_s1[22] ) );
  HS65_GS_HA1X4 U1612 ( .A0(n1494), .B0(n1493), .CO(n1492), .S0(n1521) );
  HS65_GSS_XNOR2X3 U1613 ( .A(n1521), .B(n1500), .Z(\mul_b2/fa1_s1[21] ) );
  HS65_GS_HA1X4 U1614 ( .A0(n1496), .B0(n1495), .CO(n1493), .S0(n1522) );
  HS65_GSS_XNOR2X3 U1615 ( .A(n1522), .B(n1502), .Z(\mul_b2/fa1_s1[20] ) );
  HS65_GS_HA1X4 U1616 ( .A0(n1498), .B0(n1497), .CO(n1495), .S0(n1523) );
  HS65_GSS_XNOR2X3 U1617 ( .A(n1523), .B(n1504), .Z(\mul_b2/fa1_s1[19] ) );
  HS65_GS_HA1X4 U1618 ( .A0(n1500), .B0(n1499), .CO(n1497), .S0(n1524) );
  HS65_GSS_XNOR2X3 U1619 ( .A(n1524), .B(n1506), .Z(\mul_b2/fa1_s1[18] ) );
  HS65_GS_HA1X4 U1620 ( .A0(n1502), .B0(n1501), .CO(n1499), .S0(n1525) );
  HS65_GSS_XNOR2X3 U1621 ( .A(n1525), .B(n1508), .Z(\mul_b2/fa1_s1[17] ) );
  HS65_GS_HA1X4 U1622 ( .A0(n1504), .B0(n1503), .CO(n1501), .S0(n1526) );
  HS65_GSS_XNOR2X3 U1623 ( .A(n1526), .B(n1510), .Z(\mul_b2/fa1_s1[16] ) );
  HS65_GS_HA1X4 U1624 ( .A0(n1506), .B0(n1505), .CO(n1503), .S0(n1527) );
  HS65_GSS_XNOR2X3 U1625 ( .A(n1527), .B(n1512), .Z(\mul_b2/fa1_s1[15] ) );
  HS65_GS_HA1X4 U1626 ( .A0(n1508), .B0(n1507), .CO(n1505), .S0(n1528) );
  HS65_GSS_XNOR2X3 U1627 ( .A(n1528), .B(n1514), .Z(\mul_b2/fa1_s1[14] ) );
  HS65_GS_HA1X4 U1628 ( .A0(n1510), .B0(n1509), .CO(n1507), .S0(n1529) );
  HS65_GSS_XNOR2X3 U1629 ( .A(n1529), .B(n1516), .Z(\mul_b2/fa1_s1[13] ) );
  HS65_GS_HA1X4 U1630 ( .A0(n1512), .B0(n1511), .CO(n1509), .S0(n1530) );
  HS65_GSS_XNOR2X3 U1631 ( .A(n1530), .B(n1518), .Z(\mul_b2/fa1_s1[12] ) );
  HS65_GS_HA1X4 U1632 ( .A0(n1514), .B0(n1513), .CO(n1511), .S0(n1531) );
  HS65_GSS_XNOR2X3 U1633 ( .A(n1531), .B(n1751), .Z(\mul_b2/fa1_s1[11] ) );
  HS65_GS_HA1X4 U1634 ( .A0(n1516), .B0(n1515), .CO(n1513), .S0(n1532) );
  HS65_GSS_XNOR2X3 U1635 ( .A(n1532), .B(n1742), .Z(\mul_b2/fa1_s1[10] ) );
  HS65_GS_HA1X4 U1636 ( .A0(n1518), .B0(n1517), .CO(n1515), .S0(n1533) );
  HS65_GSS_XNOR2X3 U1637 ( .A(n1533), .B(n1741), .Z(\mul_b2/fa1_s1[9] ) );
  HS65_GS_AND2X4 U1638 ( .A(x_reg2[14]), .B(n1519), .Z(\mul_b2/fa1_c1[23] ) );
  HS65_GS_AND2X4 U1639 ( .A(n1520), .B(x_reg2[13]), .Z(\mul_b2/fa1_c1[22] ) );
  HS65_GS_AND2X4 U1640 ( .A(x_reg2[12]), .B(n1521), .Z(\mul_b2/fa1_c1[21] ) );
  HS65_GS_AND2X4 U1641 ( .A(x_reg2[11]), .B(n1522), .Z(\mul_b2/fa1_c1[20] ) );
  HS65_GS_AND2X4 U1642 ( .A(x_reg2[10]), .B(n1523), .Z(\mul_b2/fa1_c1[19] ) );
  HS65_GS_AND2X4 U1643 ( .A(x_reg2[9]), .B(n1524), .Z(\mul_b2/fa1_c1[18] ) );
  HS65_GS_AND2X4 U1644 ( .A(x_reg2[8]), .B(n1525), .Z(\mul_b2/fa1_c1[17] ) );
  HS65_GS_AND2X4 U1645 ( .A(x_reg2[7]), .B(n1526), .Z(\mul_b2/fa1_c1[16] ) );
  HS65_GS_AND2X4 U1646 ( .A(x_reg2[6]), .B(n1527), .Z(\mul_b2/fa1_c1[15] ) );
  HS65_GS_AND2X4 U1647 ( .A(x_reg2[5]), .B(n1528), .Z(\mul_b2/fa1_c1[14] ) );
  HS65_GS_AND2X4 U1648 ( .A(x_reg2[4]), .B(n1529), .Z(\mul_b2/fa1_c1[13] ) );
  HS65_GS_AND2X4 U1649 ( .A(x_reg2[3]), .B(n1530), .Z(\mul_b2/fa1_c1[12] ) );
  HS65_GS_AND2X4 U1650 ( .A(x_reg2[2]), .B(n1531), .Z(\mul_b2/fa1_c1[11] ) );
  HS65_GS_AND2X4 U1651 ( .A(x_reg2[1]), .B(n1532), .Z(\mul_b2/fa1_c1[10] ) );
  HS65_GS_AND2X4 U1652 ( .A(x_reg2[0]), .B(n1533), .Z(\mul_b2/fa1_c1[9] ) );
  HS65_GS_IVX2 U1653 ( .A(n1571), .Z(n1790) );
  HS65_GS_FA1X4 U1654 ( .A0(n1536), .B0(n1535), .CI(n1534), .CO(n827), .S0(
        n1537) );
  HS65_GS_OAI21X2 U1655 ( .A(n1790), .B(n1537), .C(n1791), .Z(
        \mul_b2/result_sat[14] ) );
  HS65_GS_FA1X4 U1656 ( .A0(n1540), .B0(n1539), .CI(n1538), .CO(n817), .S0(
        n1541) );
  HS65_GS_AO12X4 U1657 ( .A(n1541), .B(n1571), .C(n1570), .Z(
        \mul_b2/result_sat[11] ) );
  HS65_GS_FA1X4 U1658 ( .A0(n1544), .B0(n1543), .CI(n1542), .CO(n1538), .S0(
        n1545) );
  HS65_GS_OA12X4 U1659 ( .A(n1570), .B(n1545), .C(n1571), .Z(
        \mul_b2/result_sat[10] ) );
  HS65_GS_FA1X4 U1660 ( .A0(n1548), .B0(n1547), .CI(n1546), .CO(n1543), .S0(
        n1549) );
  HS65_GS_AO12X4 U1661 ( .A(n1549), .B(n1571), .C(n1570), .Z(
        \mul_b2/result_sat[9] ) );
  HS65_GS_FA1X4 U1662 ( .A0(n1552), .B0(n1551), .CI(n1550), .CO(n1546), .S0(
        n1553) );
  HS65_GS_AO12X4 U1663 ( .A(n1553), .B(n1571), .C(n1570), .Z(
        \mul_b2/result_sat[8] ) );
  HS65_GSS_XOR2X3 U1664 ( .A(n1555), .B(n1554), .Z(n1556) );
  HS65_GSS_XNOR2X3 U1665 ( .A(n1557), .B(n1556), .Z(n1558) );
  HS65_GS_OAI21X2 U1666 ( .A(n1790), .B(n1558), .C(n1791), .Z(
        \mul_b2/result_sat[6] ) );
  HS65_GS_OAI21X2 U1667 ( .A(n1561), .B(n1560), .C(n1559), .Z(n1562) );
  HS65_GS_OAI21X2 U1668 ( .A(n1790), .B(n1562), .C(n1791), .Z(
        \mul_b2/result_sat[5] ) );
  HS65_GS_FA1X4 U1669 ( .A0(n1565), .B0(n1564), .CI(n1563), .CO(n356), .S0(
        n1566) );
  HS65_GS_AO12X4 U1670 ( .A(n1566), .B(n1571), .C(n1570), .Z(
        \mul_b2/result_sat[4] ) );
  HS65_GS_FA1X4 U1671 ( .A0(n1569), .B0(n1568), .CI(n1567), .CO(n1563), .S0(
        n1572) );
  HS65_GS_AO12X4 U1672 ( .A(n1572), .B(n1571), .C(n1570), .Z(
        \mul_b2/result_sat[3] ) );
  HS65_GS_OAI21X2 U1673 ( .A(n1575), .B(n1574), .C(n1573), .Z(n1576) );
  HS65_GS_OAI21X2 U1674 ( .A(n1790), .B(n1576), .C(n1791), .Z(
        \mul_b2/result_sat[1] ) );
  HS65_GS_OAI21X2 U1675 ( .A(n1579), .B(n1578), .C(n1577), .Z(n1580) );
  HS65_GS_OAI21X2 U1676 ( .A(n1790), .B(n1580), .C(n1791), .Z(
        \mul_b2/result_sat[0] ) );
  HS65_GS_AND2X4 U1677 ( .A(x_z2[14]), .B(n1581), .Z(\mul_b1/fa1_c2[28] ) );
  HS65_GS_AND2X4 U1678 ( .A(x_z2[13]), .B(n1582), .Z(\mul_b1/fa1_c2[27] ) );
  HS65_GS_AND2X4 U1679 ( .A(x_z2[12]), .B(n1583), .Z(\mul_b1/fa1_c2[26] ) );
  HS65_GS_AND2X4 U1680 ( .A(x_z2[11]), .B(n1584), .Z(\mul_b1/fa1_c2[25] ) );
  HS65_GS_AND2X4 U1681 ( .A(x_z2[10]), .B(n1585), .Z(\mul_b1/fa1_c2[24] ) );
  HS65_GS_AND2X4 U1682 ( .A(x_z2[9]), .B(n1586), .Z(\mul_b1/fa1_c2[23] ) );
  HS65_GS_AND2X4 U1683 ( .A(x_z2[8]), .B(n1587), .Z(\mul_b1/fa1_c2[22] ) );
  HS65_GS_AND2X4 U1684 ( .A(x_z2[7]), .B(n1588), .Z(\mul_b1/fa1_c2[21] ) );
  HS65_GS_AND2X4 U1685 ( .A(x_z2[6]), .B(n1589), .Z(\mul_b1/fa1_c2[20] ) );
  HS65_GS_AND2X4 U1686 ( .A(x_z2[5]), .B(n1590), .Z(\mul_b1/fa1_c2[19] ) );
  HS65_GS_AND2X4 U1687 ( .A(x_z2[4]), .B(n1591), .Z(\mul_b1/fa1_c2[18] ) );
  HS65_GS_AND2X4 U1688 ( .A(x_z2[3]), .B(n1592), .Z(\mul_b1/fa1_c2[17] ) );
  HS65_GS_AND2X4 U1689 ( .A(x_z2[2]), .B(n1593), .Z(\mul_b1/fa1_c2[16] ) );
  HS65_GS_AND2X4 U1690 ( .A(x_z2[1]), .B(n1594), .Z(\mul_b1/fa1_c2[15] ) );
  HS65_GS_AND2X4 U1691 ( .A(x_z2[0]), .B(n1595), .Z(\mul_b1/fa1_c2[14] ) );
  HS65_GS_FA1X4 U1692 ( .A0(n1598), .B0(n1597), .CI(n1596), .CO(n1604), .S0(
        n1618) );
  HS65_GS_FA1X4 U1693 ( .A0(n1601), .B0(n1600), .CI(n1599), .CO(n1013), .S0(
        n1617) );
  HS65_GS_FA1X4 U1694 ( .A0(n1604), .B0(n1603), .CI(n1602), .CO(n1609), .S0(
        n1614) );
  HS65_GS_FA1X4 U1695 ( .A0(n1607), .B0(n1606), .CI(n1605), .CO(n1600), .S0(
        n1613) );
  HS65_GS_FA1X4 U1696 ( .A0(n1610), .B0(n1609), .CI(n1608), .CO(n1606), .S0(
        n1612) );
  HS65_GS_AND3X4 U1697 ( .A(n1614), .B(n1613), .C(n1612), .Z(n1611) );
  HS65_GS_IVX2 U1698 ( .A(\mul_a1/result_sat[15] ), .Z(n1615) );
  HS65_GS_AOI12X2 U1699 ( .A(n1617), .B(n1611), .C(n1615), .Z(n1784) );
  HS65_GS_IVX2 U1700 ( .A(n1784), .Z(n1655) );
  HS65_GS_OR3X4 U1701 ( .A(n1614), .B(n1613), .C(n1612), .Z(n1616) );
  HS65_GS_OAI21X2 U1702 ( .A(n1617), .B(n1616), .C(n1615), .Z(n1785) );
  HS65_GS_IVX2 U1703 ( .A(n1785), .Z(n1646) );
  HS65_GS_AO12X4 U1704 ( .A(n1618), .B(n1655), .C(n1646), .Z(
        \mul_a1/result_sat[14] ) );
  HS65_GS_FA1X4 U1705 ( .A0(n1621), .B0(n1620), .CI(n1619), .CO(n1597), .S0(
        n1622) );
  HS65_GS_OA12X4 U1706 ( .A(n1646), .B(n1622), .C(n1655), .Z(
        \mul_a1/result_sat[13] ) );
  HS65_GS_FA1X4 U1707 ( .A0(n1625), .B0(n1624), .CI(n1623), .CO(n1620), .S0(
        n1626) );
  HS65_GS_AO12X4 U1708 ( .A(n1626), .B(n1655), .C(n1646), .Z(
        \mul_a1/result_sat[12] ) );
  HS65_GS_FA1X4 U1709 ( .A0(n1629), .B0(n1628), .CI(n1627), .CO(n1624), .S0(
        n1630) );
  HS65_GS_OA12X4 U1710 ( .A(n1646), .B(n1630), .C(n1655), .Z(
        \mul_a1/result_sat[11] ) );
  HS65_GS_FA1X4 U1711 ( .A0(n1633), .B0(n1632), .CI(n1631), .CO(n1629), .S0(
        n1634) );
  HS65_GS_AO12X4 U1712 ( .A(n1634), .B(n1655), .C(n1646), .Z(
        \mul_a1/result_sat[10] ) );
  HS65_GS_FA1X4 U1713 ( .A0(n1637), .B0(n1636), .CI(n1635), .CO(n1632), .S0(
        n1638) );
  HS65_GS_OA12X4 U1714 ( .A(n1646), .B(n1638), .C(n1655), .Z(
        \mul_a1/result_sat[9] ) );
  HS65_GS_FA1X4 U1715 ( .A0(n1641), .B0(n1640), .CI(n1639), .CO(n1637), .S0(
        n1642) );
  HS65_GS_OA12X4 U1716 ( .A(n1646), .B(n1642), .C(n1655), .Z(
        \mul_a1/result_sat[8] ) );
  HS65_GS_FA1X4 U1717 ( .A0(n1645), .B0(n1644), .CI(n1643), .CO(n1640), .S0(
        n1647) );
  HS65_GS_AO12X4 U1718 ( .A(n1647), .B(n1655), .C(n1646), .Z(
        \mul_a1/result_sat[7] ) );
  HS65_GSS_XNOR2X3 U1719 ( .A(n1649), .B(n1648), .Z(n1651) );
  HS65_GS_OAI21X2 U1720 ( .A(n1651), .B(n1652), .C(n1785), .Z(n1650) );
  HS65_GS_CB4I1X4 U1721 ( .A(n1652), .B(n1651), .C(n1650), .D(n1655), .Z(
        \mul_a1/result_sat[6] ) );
  HS65_GSS_XNOR2X3 U1722 ( .A(n1654), .B(n1653), .Z(n1657) );
  HS65_GS_OAI21X2 U1723 ( .A(n1657), .B(n1658), .C(n1785), .Z(n1656) );
  HS65_GS_CB4I1X4 U1724 ( .A(n1658), .B(n1657), .C(n1656), .D(n1655), .Z(
        \mul_a1/result_sat[5] ) );
  HS65_GSS_XOR3X2 U1725 ( .A(n1659), .B(\DP_OP_371J1_181_1383/n79 ), .C(
        x_reg2[14]), .Z(\mul_b2/fa1_s0[18] ) );
  HS65_GSS_XOR3X2 U1726 ( .A(\DP_OP_371J1_181_1383/n79 ), .B(x_reg2[13]), .C(
        n1660), .Z(\mul_b2/fa1_s0[17] ) );
  HS65_GSS_XOR3X2 U1727 ( .A(\DP_OP_371J1_181_1383/n79 ), .B(x_reg2[12]), .C(
        n1661), .Z(\mul_b2/fa1_s0[16] ) );
  HS65_GSS_XOR3X2 U1728 ( .A(\DP_OP_371J1_181_1383/n79 ), .B(x_reg2[11]), .C(
        n1662), .Z(\mul_b2/fa1_s0[15] ) );
  HS65_GSS_XOR3X2 U1729 ( .A(x_reg2[14]), .B(x_reg2[10]), .C(n1663), .Z(
        \mul_b2/fa1_s0[14] ) );
  HS65_GSS_XOR3X2 U1730 ( .A(x_reg2[13]), .B(x_reg2[9]), .C(n1664), .Z(
        \mul_b2/fa1_s0[13] ) );
  HS65_GSS_XOR3X2 U1731 ( .A(x_reg2[12]), .B(x_reg2[8]), .C(n1665), .Z(
        \mul_b2/fa1_s0[12] ) );
  HS65_GSS_XOR3X2 U1732 ( .A(x_reg2[11]), .B(x_reg2[7]), .C(n1666), .Z(
        \mul_b2/fa1_s0[11] ) );
  HS65_GSS_XOR3X2 U1733 ( .A(x_reg2[10]), .B(x_reg2[6]), .C(n1667), .Z(
        \mul_b2/fa1_s0[10] ) );
  HS65_GSS_XOR3X2 U1734 ( .A(x_reg2[9]), .B(x_reg2[5]), .C(n1668), .Z(
        \mul_b2/fa1_s0[9] ) );
  HS65_GSS_XOR3X2 U1735 ( .A(x_reg2[8]), .B(x_reg2[4]), .C(n1669), .Z(
        \mul_b2/fa1_s0[8] ) );
  HS65_GSS_XOR3X2 U1736 ( .A(x_reg2[7]), .B(x_reg2[3]), .C(n1670), .Z(
        \mul_b2/fa1_s0[7] ) );
  HS65_GSS_XOR3X2 U1737 ( .A(x_reg2[6]), .B(x_reg2[2]), .C(n1671), .Z(
        \mul_b2/fa1_s0[6] ) );
  HS65_GSS_XOR3X2 U1738 ( .A(x_reg2[5]), .B(x_reg2[1]), .C(n1672), .Z(
        \mul_b2/fa1_s0[5] ) );
  HS65_GSS_XOR3X2 U1739 ( .A(x_reg2[4]), .B(x_reg2[0]), .C(n1673), .Z(
        \mul_b2/fa1_s0[4] ) );
  HS65_GS_AND2X4 U1740 ( .A(x_z2[2]), .B(x_z2[0]), .Z(n1816) );
  HS65_GS_AND2X4 U1741 ( .A(x_z2[4]), .B(x_z2[2]), .Z(n1817) );
  HS65_GS_AND2X4 U1742 ( .A(x_z2[3]), .B(x_z2[1]), .Z(n1818) );
  HS65_GSS_XNOR2X3 U1743 ( .A(y_z2[15]), .B(n1674), .Z(\C63/DATA4_26 ) );
  HS65_GS_HA1X4 U1744 ( .A0(n1676), .B0(n1675), .CO(n1674), .S0(\C63/DATA4_25 ) );
  HS65_GS_HA1X4 U1745 ( .A0(n1678), .B0(n1677), .CO(n1675), .S0(\C63/DATA4_24 ) );
  HS65_GS_HA1X4 U1746 ( .A0(n1680), .B0(n1679), .CO(n1677), .S0(\C63/DATA4_23 ) );
  HS65_GS_HA1X4 U1747 ( .A0(n1682), .B0(n1681), .CO(n1679), .S0(\C63/DATA4_22 ) );
  HS65_GS_HA1X4 U1748 ( .A0(n1684), .B0(n1683), .CO(n1681), .S0(\C63/DATA4_21 ) );
  HS65_GS_HA1X4 U1749 ( .A0(n1686), .B0(n1685), .CO(n1683), .S0(\C63/DATA4_20 ) );
  HS65_GS_HA1X4 U1750 ( .A0(n1688), .B0(n1687), .CO(n1685), .S0(\C63/DATA4_19 ) );
  HS65_GS_HA1X4 U1751 ( .A0(n1690), .B0(n1689), .CO(n1687), .S0(\C63/DATA4_18 ) );
  HS65_GS_HA1X4 U1752 ( .A0(n1692), .B0(n1691), .CO(n1689), .S0(\C63/DATA4_17 ) );
  HS65_GS_HA1X4 U1753 ( .A0(n1694), .B0(n1693), .CO(n1691), .S0(\C63/DATA4_16 ) );
  HS65_GS_HA1X4 U1754 ( .A0(n1696), .B0(n1695), .CO(n1693), .S0(\C63/DATA4_15 ) );
  HS65_GS_HA1X4 U1755 ( .A0(n1698), .B0(n1697), .CO(n1695), .S0(\C63/DATA4_14 ) );
  HS65_GS_HA1X4 U1756 ( .A0(n1700), .B0(n1699), .CO(n1697), .S0(\C63/DATA4_13 ) );
  HS65_GS_HA1X4 U1757 ( .A0(n1702), .B0(n1701), .CO(n1699), .S0(\C63/DATA4_12 ) );
  HS65_GSS_XNOR2X3 U1758 ( .A(y_z1[15]), .B(n1703), .Z(\C56/DATA4_30 ) );
  HS65_GS_HA1X4 U1759 ( .A0(n1705), .B0(n1704), .CO(n1703), .S0(\C56/DATA4_29 ) );
  HS65_GS_HA1X4 U1760 ( .A0(n1724), .B0(n1706), .CO(n1704), .S0(\C56/DATA4_28 ) );
  HS65_GS_HA1X4 U1761 ( .A0(n1726), .B0(n1707), .CO(n1706), .S0(\C56/DATA4_27 ) );
  HS65_GS_HA1X4 U1762 ( .A0(n1728), .B0(n1708), .CO(n1707), .S0(\C56/DATA4_26 ) );
  HS65_GS_HA1X4 U1763 ( .A0(n1730), .B0(n1709), .CO(n1708), .S0(\C56/DATA4_25 ) );
  HS65_GS_HA1X4 U1764 ( .A0(n1732), .B0(n1710), .CO(n1709), .S0(\C56/DATA4_24 ) );
  HS65_GS_HA1X4 U1765 ( .A0(n1734), .B0(n1711), .CO(n1710), .S0(\C56/DATA4_23 ) );
  HS65_GS_HA1X4 U1766 ( .A0(n1736), .B0(n1712), .CO(n1711), .S0(\C56/DATA4_22 ) );
  HS65_GS_HA1X4 U1767 ( .A0(n1738), .B0(n1713), .CO(n1712), .S0(\C56/DATA4_21 ) );
  HS65_GS_HA1X4 U1768 ( .A0(n1740), .B0(n1714), .CO(n1713), .S0(\C56/DATA4_20 ) );
  HS65_GS_HA1X4 U1769 ( .A0(n1716), .B0(n1715), .CO(n1714), .S0(\C56/DATA4_19 ) );
  HS65_GS_HA1X4 U1770 ( .A0(n1718), .B0(n1717), .CO(n1715), .S0(\C56/DATA4_18 ) );
  HS65_GS_HA1X4 U1771 ( .A0(n1720), .B0(n1719), .CO(n1717), .S0(\C56/DATA4_17 ) );
  HS65_GS_HA1X4 U1772 ( .A0(n1754), .B0(n1721), .CO(n1719), .S0(\C56/DATA4_16 ) );
  HS65_GS_HA1X4 U1773 ( .A0(n1755), .B0(n1753), .CO(n1721), .S0(\C56/DATA4_15 ) );
  HS65_GSS_XNOR2X3 U1774 ( .A(y_z1[15]), .B(n1722), .Z(\C49/DATA3_16 ) );
  HS65_GS_HA1X4 U1775 ( .A0(n1724), .B0(n1723), .CO(n1722), .S0(\C49/DATA3_15 ) );
  HS65_GS_HA1X4 U1776 ( .A0(n1726), .B0(n1725), .CO(n1723), .S0(\C49/DATA3_14 ) );
  HS65_GS_HA1X4 U1777 ( .A0(n1728), .B0(n1727), .CO(n1725), .S0(\C49/DATA3_13 ) );
  HS65_GS_HA1X4 U1778 ( .A0(n1730), .B0(n1729), .CO(n1727), .S0(\C49/DATA3_12 ) );
  HS65_GS_HA1X4 U1779 ( .A0(n1732), .B0(n1731), .CO(n1729), .S0(\C49/DATA3_11 ) );
  HS65_GS_HA1X4 U1780 ( .A0(n1734), .B0(n1733), .CO(n1731), .S0(\C49/DATA3_10 ) );
  HS65_GS_HA1X4 U1781 ( .A0(n1736), .B0(n1735), .CO(n1733), .S0(\C49/DATA3_9 )
         );
  HS65_GS_HA1X4 U1782 ( .A0(n1738), .B0(n1737), .CO(n1735), .S0(\C49/DATA3_8 )
         );
  HS65_GS_HA1X4 U1783 ( .A0(n1740), .B0(n1739), .CO(n1737), .S0(\C49/DATA3_7 )
         );
  HS65_GS_HA1X4 U1784 ( .A0(n1742), .B0(n1741), .CO(n1750), .S0(
        \mul_b2/fa1_s1[7] ) );
  HS65_GSS_XNOR2X3 U1785 ( .A(\DP_OP_331J1_157_5454/n87 ), .B(n1743), .Z(
        \C33/DATA4_20 ) );
  HS65_GS_HA1X4 U1786 ( .A0(n1745), .B0(n1744), .CO(n1743), .S0(\C33/DATA4_19 ) );
  HS65_GS_HA1X4 U1787 ( .A0(n1747), .B0(n1746), .CO(n1744), .S0(\C33/DATA4_18 ) );
  HS65_GS_HA1X4 U1788 ( .A0(n1749), .B0(n1748), .CO(n1746), .S0(\C33/DATA4_17 ) );
  HS65_GS_HA1X4 U1789 ( .A0(n1751), .B0(n1750), .CO(n1517), .S0(\C43/DATA4_8 )
         );
  HS65_GS_HA1X4 U1790 ( .A0(n1752), .B0(n1411), .CO(n1252), .S0(
        \mul_b1/fa1_s1[7] ) );
  HS65_GS_AOI12X2 U1791 ( .A(n1753), .B(n1755), .C(\mul_a1/fa1_c1[8] ), .Z(
        \mul_a1/fa1_s1[8] ) );
  HS65_GS_AOI12X2 U1792 ( .A(n1755), .B(n1754), .C(\mul_a1/fa1_c1[9] ), .Z(
        \mul_a1/fa1_s1[9] ) );
  HS65_GS_FA1X4 U1793 ( .A0(\mul_a1/fa1_s1[7] ), .B0(y_z1[3]), .CI(y_z1[2]), 
        .CO(\mul_a1/fa1_c1[10] ), .S0(\mul_a1/fa1_s1[10] ) );
  HS65_GS_FA1X4 U1794 ( .A0(y_z1[4]), .B0(y_z1[3]), .CI(y_z1[1]), .CO(
        \mul_a1/fa1_c1[11] ), .S0(\mul_a1/fa1_s1[11] ) );
  HS65_GS_FA1X4 U1795 ( .A0(y_z1[5]), .B0(y_z1[4]), .CI(y_z1[2]), .CO(
        \mul_a1/fa1_c1[12] ), .S0(\mul_a1/fa1_s1[12] ) );
  HS65_GS_FA1X4 U1796 ( .A0(y_z1[6]), .B0(y_z1[5]), .CI(y_z1[3]), .CO(
        \mul_a1/fa1_c1[13] ), .S0(\mul_a1/fa1_s1[13] ) );
  HS65_GS_FA1X4 U1797 ( .A0(y_z1[7]), .B0(y_z1[6]), .CI(y_z1[4]), .CO(
        \mul_a1/fa1_c1[14] ), .S0(\mul_a1/fa1_s1[14] ) );
  HS65_GS_FA1X4 U1798 ( .A0(y_z1[8]), .B0(y_z1[7]), .CI(y_z1[5]), .CO(
        \mul_a1/fa1_c1[15] ), .S0(\mul_a1/fa1_s1[15] ) );
  HS65_GS_FA1X4 U1799 ( .A0(y_z1[9]), .B0(y_z1[8]), .CI(y_z1[6]), .CO(
        \mul_a1/fa1_c1[16] ), .S0(\mul_a1/fa1_s1[16] ) );
  HS65_GS_FA1X4 U1800 ( .A0(y_z1[10]), .B0(y_z1[9]), .CI(y_z1[7]), .CO(
        \mul_a1/fa1_c1[17] ), .S0(\mul_a1/fa1_s1[17] ) );
  HS65_GS_FA1X4 U1801 ( .A0(y_z1[11]), .B0(y_z1[10]), .CI(y_z1[8]), .CO(
        \mul_a1/fa1_c1[18] ), .S0(\mul_a1/fa1_s1[18] ) );
  HS65_GS_FA1X4 U1802 ( .A0(y_z1[12]), .B0(y_z1[11]), .CI(y_z1[9]), .CO(
        \mul_a1/fa1_c1[19] ), .S0(\mul_a1/fa1_s1[19] ) );
  HS65_GS_FA1X4 U1803 ( .A0(y_z1[13]), .B0(y_z1[12]), .CI(y_z1[10]), .CO(
        \mul_a1/fa1_c1[20] ), .S0(\mul_a1/fa1_s1[20] ) );
  HS65_GS_FA1X4 U1804 ( .A0(y_z1[14]), .B0(y_z1[13]), .CI(y_z1[11]), .CO(
        \mul_a1/fa1_c1[21] ), .S0(\mul_a1/fa1_s1[21] ) );
  HS65_GS_FA1X4 U1805 ( .A0(y_z1[15]), .B0(y_z1[14]), .CI(y_z1[12]), .CO(
        \mul_a1/fa1_c1[22] ), .S0(\mul_a1/fa1_s1[22] ) );
  HS65_GS_IVX2 U1806 ( .A(n1756), .Z(n1761) );
  HS65_GS_IVX2 U1807 ( .A(n1757), .Z(n1759) );
  HS65_GS_AOI22X1 U1808 ( .A(n1761), .B(n1760), .C(n1759), .D(n1758), .Z(n1764) );
  HS65_GS_AOI12X2 U1809 ( .A(n1764), .B(n1763), .C(n1762), .Z(
        \mul_a2/result_sat[1] ) );
  HS65_GS_AOI12X2 U1810 ( .A(n1767), .B(n1766), .C(n1765), .Z(n1768) );
  HS65_GS_AOI12X2 U1811 ( .A(n1768), .B(n1785), .C(n1784), .Z(
        \mul_a1/result_sat[0] ) );
  HS65_GS_AOI12X2 U1812 ( .A(n1771), .B(n1770), .C(n1769), .Z(n1772) );
  HS65_GS_AOI12X2 U1813 ( .A(n1772), .B(n1785), .C(n1784), .Z(
        \mul_a1/result_sat[1] ) );
  HS65_GS_AOI12X2 U1814 ( .A(n1775), .B(n1774), .C(n1773), .Z(n1776) );
  HS65_GS_AOI12X2 U1815 ( .A(n1776), .B(n1785), .C(n1784), .Z(
        \mul_a1/result_sat[2] ) );
  HS65_GS_AOI12X2 U1816 ( .A(n1779), .B(n1778), .C(n1777), .Z(n1780) );
  HS65_GS_AOI12X2 U1817 ( .A(n1780), .B(n1785), .C(n1784), .Z(
        \mul_a1/result_sat[3] ) );
  HS65_GS_AOI12X2 U1818 ( .A(n1783), .B(n1782), .C(n1781), .Z(n1786) );
  HS65_GS_AOI12X2 U1819 ( .A(n1786), .B(n1785), .C(n1784), .Z(
        \mul_a1/result_sat[4] ) );
  HS65_GS_FA1X4 U1820 ( .A0(n1789), .B0(n1788), .CI(n1787), .CO(n1535), .S0(
        n1792) );
  HS65_GS_AOI12X2 U1821 ( .A(n1792), .B(n1791), .C(n1790), .Z(
        \mul_b2/result_sat[13] ) );
  HS65_GS_FA1X4 U1822 ( .A0(n1795), .B0(n1794), .CI(n1793), .CO(n515), .S0(
        n1798) );
  HS65_GS_AOI12X2 U1823 ( .A(n1798), .B(n1797), .C(n1796), .Z(
        \mul_b1/result_sat[0] ) );
  HS65_GS_IVX2 U1824 ( .A(n1799), .Z(n1804) );
  HS65_GS_IVX2 U1825 ( .A(n1800), .Z(n1802) );
  HS65_GS_AOI22X1 U1826 ( .A(n1804), .B(n1803), .C(n1802), .D(n1801), .Z(n1807) );
  HS65_GS_AOI12X2 U1827 ( .A(n1807), .B(n1806), .C(n1805), .Z(
        \mul_b0/result_sat[1] ) );
  HS65_GS_AOI12X2 U1828 ( .A(n1810), .B(n1809), .C(n1808), .Z(n1870) );
endmodule


module opti_sos_3 ( clk, rst_n, data_in, valid_in, b0, b1, b2, a1, a2, 
        data_out, valid_out );
  input [15:0] data_in;
  input [15:0] b0;
  input [15:0] b1;
  input [15:0] b2;
  input [15:0] a1;
  input [15:0] a2;
  output [15:0] data_out;
  input clk, rst_n, valid_in;
  output valid_out;
  wire   valid_T1, valid_T3, valid_T2, \mul_b0/result_sat[15] ,
         \mul_b0/result_sat[14] , \mul_b0/result_sat[13] ,
         \mul_b0/result_sat[12] , \mul_b0/result_sat[11] ,
         \mul_b0/result_sat[10] , \mul_b0/result_sat[9] ,
         \mul_b0/result_sat[8] , \mul_b0/result_sat[7] ,
         \mul_b0/result_sat[6] , \mul_b0/result_sat[5] ,
         \mul_b0/result_sat[4] , \mul_b0/result_sat[3] ,
         \mul_b0/result_sat[2] , \mul_b0/result_sat[1] ,
         \mul_b0/result_sat[0] , \mul_b0/fa1_s2_r[33] , \mul_b0/fa1_s2_r[32] ,
         \mul_b0/fa1_s2_r[31] , \mul_b0/fa1_s2_r[30] , \mul_b0/fa1_s2_r[29] ,
         \mul_b0/fa1_s2_r[28] , \mul_b0/fa1_s2_r[27] , \mul_b0/fa1_s2_r[26] ,
         \mul_b0/fa1_s2_r[25] , \mul_b0/fa1_s2_r[24] , \mul_b0/fa1_s2_r[23] ,
         \mul_b0/fa1_s2_r[22] , \mul_b0/fa1_s2_r[21] , \mul_b0/fa1_s2_r[20] ,
         \mul_b0/fa1_s2_r[19] , \mul_b0/fa1_s2_r[18] , \mul_b0/fa1_s2_r[17] ,
         \mul_b0/fa1_s2_r[16] , \mul_b0/fa1_s2_r[15] , \mul_b0/fa1_s2_r[14] ,
         \mul_b0/fa1_s2_r[13] , \mul_b0/fa1_s2_r[12] , \mul_b0/fa1_s1_r[33] ,
         \mul_b0/fa1_s1_r[32] , \mul_b0/fa1_s1_r[31] , \mul_b0/fa1_s1_r[30] ,
         \mul_b0/fa1_s1_r[29] , \mul_b0/fa1_s1_r[28] , \mul_b0/fa1_s1_r[27] ,
         \mul_b0/fa1_s1_r[26] , \mul_b0/fa1_s1_r[25] , \mul_b0/fa1_s1_r[24] ,
         \mul_b0/fa1_s1_r[23] , \mul_b0/fa1_s1_r[22] , \mul_b0/fa1_s1_r[21] ,
         \mul_b0/fa1_s1_r[20] , \mul_b0/fa1_s1_r[19] , \mul_b0/fa1_s1_r[18] ,
         \mul_b0/fa1_s1_r[17] , \mul_b0/fa1_s1_r[16] , \mul_b0/fa1_s1_r[15] ,
         \mul_b0/fa1_s1_r[14] , \mul_b0/fa1_s1_r[13] , \mul_b0/fa1_s1_r[12] ,
         \mul_b0/fa1_s1_r[11] , \mul_b0/fa1_s1_r[10] , \mul_b0/fa1_s1_r[9] ,
         \mul_b0/fa1_s1_r[8] , \mul_b0/fa1_c0_r[20] , \mul_b0/fa1_c0_r[19] ,
         \mul_b0/fa1_c0_r[18] , \mul_b0/fa1_c0_r[17] , \mul_b0/fa1_c0_r[16] ,
         \mul_b0/fa1_c0_r[15] , \mul_b0/fa1_c0_r[14] , \mul_b0/fa1_c0_r[13] ,
         \mul_b0/fa1_c0_r[12] , \mul_b0/fa1_c0_r[11] , \mul_b0/fa1_c0_r[10] ,
         \mul_b0/fa1_c0_r[9] , \mul_b0/fa1_c0_r[8] , \mul_b0/fa1_c0_r[7] ,
         \mul_b0/fa1_c0_r[6] , \mul_b0/fa1_c0_r[5] , \mul_b0/fa1_s0_r[33] ,
         \mul_b0/fa1_s0_r[32] , \mul_b0/fa1_s0_r[31] , \mul_b0/fa1_s0_r[30] ,
         \mul_b0/fa1_s0_r[29] , \mul_b0/fa1_s0_r[28] , \mul_b0/fa1_s0_r[27] ,
         \mul_b0/fa1_s0_r[26] , \mul_b0/fa1_s0_r[25] , \mul_b0/fa1_s0_r[24] ,
         \mul_b0/fa1_s0_r[23] , \mul_b0/fa1_s0_r[22] , \mul_b0/fa1_s0_r[21] ,
         \mul_b0/fa1_s0_r[20] , \mul_b0/fa1_s0_r[19] , \mul_b0/fa1_s0_r[18] ,
         \mul_b0/fa1_s0_r[17] , \mul_b0/fa1_s0_r[16] , \mul_b0/fa1_s0_r[15] ,
         \mul_b0/fa1_s0_r[14] , \mul_b0/fa1_s0_r[13] , \mul_b0/fa1_s0_r[12] ,
         \mul_b0/fa1_s0_r[11] , \mul_b0/fa1_s0_r[10] , \mul_b0/fa1_s0_r[9] ,
         \mul_b0/fa1_s0_r[8] , \mul_b0/fa1_s0_r[7] , \mul_b0/fa1_s0_r[6] ,
         \mul_b0/fa1_c0[20] , \mul_b0/fa1_c0[19] , \mul_b0/fa1_c0[18] ,
         \mul_b0/fa1_c0[17] , \mul_b0/fa1_c0[16] , \mul_b0/fa1_c0[15] ,
         \mul_b0/fa1_c0[14] , \mul_b0/fa1_c0[13] , \mul_b0/fa1_c0[12] ,
         \mul_b0/fa1_c0[11] , \mul_b0/fa1_c0[10] , \mul_b0/fa1_c0[9] ,
         \mul_b0/fa1_c0[8] , \mul_b0/fa1_c0[7] , \mul_b0/fa1_c0[6] ,
         \mul_b0/fa1_c0[5] , \mul_b0/fa1_s0[31] , \mul_b0/fa1_s0[20] ,
         \mul_b0/fa1_s0[19] , \mul_b0/fa1_s0[18] , \mul_b0/fa1_s0[17] ,
         \mul_b0/fa1_s0[16] , \mul_b0/fa1_s0[15] , \mul_b0/fa1_s0[14] ,
         \mul_b0/fa1_s0[13] , \mul_b0/fa1_s0[12] , \mul_b0/fa1_s0[11] ,
         \mul_b0/fa1_s0[10] , \mul_b0/fa1_s0[9] , \mul_b0/fa1_s0[8] ,
         \mul_b0/fa1_s0[7] , \mul_b0/fa1_s0[6] , \mul_b1/result_sat[15] ,
         \mul_b1/result_sat[14] , \mul_b1/result_sat[13] ,
         \mul_b1/result_sat[12] , \mul_b1/result_sat[11] ,
         \mul_b1/result_sat[10] , \mul_b1/result_sat[9] ,
         \mul_b1/result_sat[8] , \mul_b1/result_sat[7] ,
         \mul_b1/result_sat[6] , \mul_b1/result_sat[5] ,
         \mul_b1/result_sat[4] , \mul_b1/result_sat[3] ,
         \mul_b1/result_sat[2] , \mul_b1/result_sat[1] ,
         \mul_b1/result_sat[0] , \mul_b1/fa1_c2_r[28] , \mul_b1/fa1_c2_r[27] ,
         \mul_b1/fa1_c2_r[26] , \mul_b1/fa1_c2_r[25] , \mul_b1/fa1_c2_r[24] ,
         \mul_b1/fa1_c2_r[23] , \mul_b1/fa1_c2_r[22] , \mul_b1/fa1_c2_r[21] ,
         \mul_b1/fa1_c2_r[20] , \mul_b1/fa1_c2_r[19] , \mul_b1/fa1_c2_r[18] ,
         \mul_b1/fa1_c2_r[17] , \mul_b1/fa1_c2_r[16] , \mul_b1/fa1_c2_r[15] ,
         \mul_b1/fa1_c2_r[14] , \mul_b1/fa1_s2_r[33] , \mul_b1/fa1_s2_r[32] ,
         \mul_b1/fa1_s2_r[31] , \mul_b1/fa1_s2_r[30] , \mul_b1/fa1_s2_r[29] ,
         \mul_b1/fa1_s2_r[28] , \mul_b1/fa1_s2_r[27] , \mul_b1/fa1_s2_r[26] ,
         \mul_b1/fa1_s2_r[25] , \mul_b1/fa1_s2_r[24] , \mul_b1/fa1_s2_r[23] ,
         \mul_b1/fa1_s2_r[22] , \mul_b1/fa1_s2_r[21] , \mul_b1/fa1_s2_r[20] ,
         \mul_b1/fa1_s2_r[19] , \mul_b1/fa1_s2_r[18] , \mul_b1/fa1_s2_r[17] ,
         \mul_b1/fa1_s2_r[16] , \mul_b1/fa1_s2_r[15] , \mul_b1/fa1_s2_r[14] ,
         \mul_b1/fa1_s2_r[13] , \mul_b1/fa1_s1_r[33] , \mul_b1/fa1_s1_r[32] ,
         \mul_b1/fa1_s1_r[31] , \mul_b1/fa1_s1_r[30] , \mul_b1/fa1_s1_r[29] ,
         \mul_b1/fa1_s1_r[28] , \mul_b1/fa1_s1_r[27] , \mul_b1/fa1_s1_r[26] ,
         \mul_b1/fa1_s1_r[25] , \mul_b1/fa1_s1_r[24] , \mul_b1/fa1_s1_r[23] ,
         \mul_b1/fa1_s1_r[22] , \mul_b1/fa1_s1_r[21] , \mul_b1/fa1_s1_r[20] ,
         \mul_b1/fa1_s1_r[19] , \mul_b1/fa1_s1_r[18] , \mul_b1/fa1_s1_r[17] ,
         \mul_b1/fa1_s1_r[16] , \mul_b1/fa1_s1_r[15] , \mul_b1/fa1_s1_r[14] ,
         \mul_b1/fa1_s1_r[13] , \mul_b1/fa1_s1_r[12] , \mul_b1/fa1_s1_r[11] ,
         \mul_b1/fa1_s1_r[10] , \mul_b1/fa1_s1_r[9] , \mul_b1/fa1_c0_r[19] ,
         \mul_b1/fa1_c0_r[18] , \mul_b1/fa1_c0_r[17] , \mul_b1/fa1_c0_r[16] ,
         \mul_b1/fa1_c0_r[15] , \mul_b1/fa1_c0_r[14] , \mul_b1/fa1_c0_r[13] ,
         \mul_b1/fa1_c0_r[12] , \mul_b1/fa1_c0_r[11] , \mul_b1/fa1_c0_r[10] ,
         \mul_b1/fa1_c0_r[9] , \mul_b1/fa1_c0_r[8] , \mul_b1/fa1_c0_r[7] ,
         \mul_b1/fa1_c0_r[6] , \mul_b1/fa1_c0_r[5] , \mul_b1/fa1_c0_r[4] ,
         \mul_b1/fa1_s0_r[33] , \mul_b1/fa1_s0_r[32] , \mul_b1/fa1_s0_r[31] ,
         \mul_b1/fa1_s0_r[30] , \mul_b1/fa1_s0_r[29] , \mul_b1/fa1_s0_r[28] ,
         \mul_b1/fa1_s0_r[27] , \mul_b1/fa1_s0_r[26] , \mul_b1/fa1_s0_r[25] ,
         \mul_b1/fa1_s0_r[24] , \mul_b1/fa1_s0_r[23] , \mul_b1/fa1_s0_r[22] ,
         \mul_b1/fa1_s0_r[21] , \mul_b1/fa1_s0_r[20] , \mul_b1/fa1_s0_r[19] ,
         \mul_b1/fa1_s0_r[18] , \mul_b1/fa1_s0_r[17] , \mul_b1/fa1_s0_r[16] ,
         \mul_b1/fa1_s0_r[15] , \mul_b1/fa1_s0_r[14] , \mul_b1/fa1_s0_r[13] ,
         \mul_b1/fa1_s0_r[12] , \mul_b1/fa1_s0_r[11] , \mul_b1/fa1_s0_r[10] ,
         \mul_b1/fa1_s0_r[9] , \mul_b1/fa1_s0_r[8] , \mul_b1/fa1_s0_r[7] ,
         \mul_b1/fa1_s0_r[6] , \mul_b1/fa1_s0_r[5] , \mul_b1/fa1_c2[28] ,
         \mul_b1/fa1_c2[27] , \mul_b1/fa1_c2[26] , \mul_b1/fa1_c2[25] ,
         \mul_b1/fa1_c2[24] , \mul_b1/fa1_c2[23] , \mul_b1/fa1_c2[22] ,
         \mul_b1/fa1_c2[21] , \mul_b1/fa1_c2[20] , \mul_b1/fa1_c2[19] ,
         \mul_b1/fa1_c2[18] , \mul_b1/fa1_c2[17] , \mul_b1/fa1_c2[16] ,
         \mul_b1/fa1_c2[15] , \mul_b1/fa1_c2[14] , \mul_b1/fa1_s2[29] ,
         \mul_b1/fa1_s2[28] , \mul_b1/fa1_s2[27] , \mul_b1/fa1_s2[26] ,
         \mul_b1/fa1_s2[25] , \mul_b1/fa1_s2[24] , \mul_b1/fa1_s2[23] ,
         \mul_b1/fa1_s2[22] , \mul_b1/fa1_s2[21] , \mul_b1/fa1_s2[20] ,
         \mul_b1/fa1_s2[19] , \mul_b1/fa1_s2[18] , \mul_b1/fa1_s2[17] ,
         \mul_b1/fa1_s2[16] , \mul_b1/fa1_s2[15] , \mul_b1/fa1_s2[14] ,
         \mul_b1/fa1_c0[19] , \mul_b1/fa1_c0[18] , \mul_b1/fa1_c0[17] ,
         \mul_b1/fa1_c0[16] , \mul_b1/fa1_c0[15] , \mul_b1/fa1_c0[14] ,
         \mul_b1/fa1_c0[13] , \mul_b1/fa1_c0[12] , \mul_b1/fa1_c0[11] ,
         \mul_b1/fa1_c0[10] , \mul_b1/fa1_c0[9] , \mul_b1/fa1_c0[8] ,
         \mul_b1/fa1_c0[7] , \mul_b1/fa1_c0[6] , \mul_b1/fa1_c0[5] ,
         \mul_b1/fa1_c0[4] , \mul_b1/fa1_s0[27] , \mul_b1/fa1_s0[20] ,
         \mul_b1/fa1_s0[19] , \mul_b1/fa1_s0[18] , \mul_b1/fa1_s0[17] ,
         \mul_b1/fa1_s0[16] , \mul_b1/fa1_s0[15] , \mul_b1/fa1_s0[14] ,
         \mul_b1/fa1_s0[13] , \mul_b1/fa1_s0[12] , \mul_b1/fa1_s0[11] ,
         \mul_b1/fa1_s0[10] , \mul_b1/fa1_s0[9] , \mul_b1/fa1_s0[8] ,
         \mul_b1/fa1_s0[7] , \mul_b1/fa1_s0[6] , \mul_b1/fa1_s0[5] ,
         \mul_b2/result_sat[15] , \mul_b2/result_sat[14] ,
         \mul_b2/result_sat[13] , \mul_b2/result_sat[12] ,
         \mul_b2/result_sat[11] , \mul_b2/result_sat[10] ,
         \mul_b2/result_sat[9] , \mul_b2/result_sat[8] ,
         \mul_b2/result_sat[7] , \mul_b2/result_sat[6] ,
         \mul_b2/result_sat[5] , \mul_b2/result_sat[4] ,
         \mul_b2/result_sat[3] , \mul_b2/result_sat[2] ,
         \mul_b2/result_sat[1] , \mul_b2/result_sat[0] , \mul_b2/fa1_s2_r[33] ,
         \mul_b2/fa1_s2_r[32] , \mul_b2/fa1_s2_r[31] , \mul_b2/fa1_s2_r[30] ,
         \mul_b2/fa1_s2_r[29] , \mul_b2/fa1_s2_r[28] , \mul_b2/fa1_s2_r[27] ,
         \mul_b2/fa1_s2_r[26] , \mul_b2/fa1_s2_r[25] , \mul_b2/fa1_s2_r[24] ,
         \mul_b2/fa1_s2_r[23] , \mul_b2/fa1_s2_r[22] , \mul_b2/fa1_s2_r[21] ,
         \mul_b2/fa1_s2_r[20] , \mul_b2/fa1_s2_r[19] , \mul_b2/fa1_s2_r[18] ,
         \mul_b2/fa1_s2_r[17] , \mul_b2/fa1_s2_r[16] , \mul_b2/fa1_s2_r[15] ,
         \mul_b2/fa1_s2_r[14] , \mul_b2/fa1_s2_r[13] , \mul_b2/fa1_s2_r[12] ,
         \mul_b2/fa1_s1_r[33] , \mul_b2/fa1_s1_r[32] , \mul_b2/fa1_s1_r[31] ,
         \mul_b2/fa1_s1_r[30] , \mul_b2/fa1_s1_r[29] , \mul_b2/fa1_s1_r[28] ,
         \mul_b2/fa1_s1_r[27] , \mul_b2/fa1_s1_r[26] , \mul_b2/fa1_s1_r[25] ,
         \mul_b2/fa1_s1_r[24] , \mul_b2/fa1_s1_r[23] , \mul_b2/fa1_s1_r[22] ,
         \mul_b2/fa1_s1_r[21] , \mul_b2/fa1_s1_r[20] , \mul_b2/fa1_s1_r[19] ,
         \mul_b2/fa1_s1_r[18] , \mul_b2/fa1_s1_r[17] , \mul_b2/fa1_s1_r[16] ,
         \mul_b2/fa1_s1_r[15] , \mul_b2/fa1_s1_r[14] , \mul_b2/fa1_s1_r[13] ,
         \mul_b2/fa1_s1_r[12] , \mul_b2/fa1_s1_r[11] , \mul_b2/fa1_s1_r[10] ,
         \mul_b2/fa1_s1_r[9] , \mul_b2/fa1_s1_r[8] , \mul_b2/fa1_c0_r[32] ,
         \mul_b2/fa1_c0_r[31] , \mul_b2/fa1_c0_r[30] , \mul_b2/fa1_c0_r[29] ,
         \mul_b2/fa1_c0_r[28] , \mul_b2/fa1_c0_r[27] , \mul_b2/fa1_c0_r[26] ,
         \mul_b2/fa1_c0_r[25] , \mul_b2/fa1_c0_r[24] , \mul_b2/fa1_c0_r[23] ,
         \mul_b2/fa1_c0_r[22] , \mul_b2/fa1_c0_r[21] , \mul_b2/fa1_c0_r[20] ,
         \mul_b2/fa1_c0_r[19] , \mul_b2/fa1_c0_r[18] , \mul_b2/fa1_c0_r[17] ,
         \mul_b2/fa1_c0_r[16] , \mul_b2/fa1_c0_r[15] , \mul_b2/fa1_c0_r[14] ,
         \mul_b2/fa1_c0_r[13] , \mul_b2/fa1_c0_r[12] , \mul_b2/fa1_c0_r[11] ,
         \mul_b2/fa1_c0_r[10] , \mul_b2/fa1_c0_r[9] , \mul_b2/fa1_c0_r[8] ,
         \mul_b2/fa1_c0_r[7] , \mul_b2/fa1_c0_r[6] , \mul_b2/fa1_c0_r[5] ,
         \mul_b2/fa1_c0_r[4] , \mul_b2/fa1_c0_r[3] , \mul_b2/fa1_c0_r[2] ,
         \mul_b2/fa1_s0_r[33] , \mul_b2/fa1_s0_r[32] , \mul_b2/fa1_s0_r[31] ,
         \mul_b2/fa1_s0_r[30] , \mul_b2/fa1_s0_r[29] , \mul_b2/fa1_s0_r[28] ,
         \mul_b2/fa1_s0_r[27] , \mul_b2/fa1_s0_r[26] , \mul_b2/fa1_s0_r[25] ,
         \mul_b2/fa1_s0_r[24] , \mul_b2/fa1_s0_r[23] , \mul_b2/fa1_s0_r[22] ,
         \mul_b2/fa1_s0_r[21] , \mul_b2/fa1_s0_r[20] , \mul_b2/fa1_s0_r[19] ,
         \mul_b2/fa1_s0_r[18] , \mul_b2/fa1_s0_r[17] , \mul_b2/fa1_s0_r[16] ,
         \mul_b2/fa1_s0_r[15] , \mul_b2/fa1_s0_r[14] , \mul_b2/fa1_s0_r[13] ,
         \mul_b2/fa1_s0_r[12] , \mul_b2/fa1_s0_r[11] , \mul_b2/fa1_s0_r[10] ,
         \mul_b2/fa1_s0_r[9] , \mul_b2/fa1_s0_r[8] , \mul_b2/fa1_s0_r[7] ,
         \mul_b2/fa1_s0_r[6] , \mul_b2/fa1_s0_r[5] , \mul_b2/fa1_s0_r[4] ,
         \mul_b2/fa1_s0_r[3] , \mul_b2/fa1_c0[16] , \mul_b2/fa1_c0[15] ,
         \mul_b2/fa1_c0[14] , \mul_b2/fa1_c0[13] , \mul_b2/fa1_c0[12] ,
         \mul_b2/fa1_c0[11] , \mul_b2/fa1_c0[10] , \mul_b2/fa1_c0[9] ,
         \mul_b2/fa1_c0[8] , \mul_b2/fa1_c0[7] , \mul_b2/fa1_c0[6] ,
         \mul_b2/fa1_c0[5] , \mul_b2/fa1_c0[4] , \mul_b2/fa1_c0[3] ,
         \mul_b2/fa1_c0[2] , \mul_b2/fa1_s0[16] , \mul_b2/fa1_s0[15] ,
         \mul_b2/fa1_s0[14] , \mul_b2/fa1_s0[13] , \mul_b2/fa1_s0[12] ,
         \mul_b2/fa1_s0[11] , \mul_b2/fa1_s0[10] , \mul_b2/fa1_s0[9] ,
         \mul_b2/fa1_s0[8] , \mul_b2/fa1_s0[7] , \mul_b2/fa1_s0[6] ,
         \mul_b2/fa1_s0[5] , \mul_b2/fa1_s0[4] , \mul_b2/fa1_s0[3] ,
         \mul_a1/result_sat[15] , \mul_a1/result_sat[14] ,
         \mul_a1/result_sat[13] , \mul_a1/result_sat[12] ,
         \mul_a1/result_sat[11] , \mul_a1/result_sat[10] ,
         \mul_a1/result_sat[9] , \mul_a1/result_sat[8] ,
         \mul_a1/result_sat[7] , \mul_a1/result_sat[6] ,
         \mul_a1/result_sat[5] , \mul_a1/result_sat[4] ,
         \mul_a1/result_sat[3] , \mul_a1/result_sat[2] ,
         \mul_a1/result_sat[1] , \mul_a1/result_sat[0] , \mul_a1/fa1_c2_r[29] ,
         \mul_a1/fa1_c2_r[28] , \mul_a1/fa1_c2_r[27] , \mul_a1/fa1_c2_r[26] ,
         \mul_a1/fa1_c2_r[25] , \mul_a1/fa1_c2_r[24] , \mul_a1/fa1_c2_r[23] ,
         \mul_a1/fa1_c2_r[22] , \mul_a1/fa1_c2_r[21] , \mul_a1/fa1_c2_r[20] ,
         \mul_a1/fa1_c2_r[19] , \mul_a1/fa1_c2_r[18] , \mul_a1/fa1_c2_r[17] ,
         \mul_a1/fa1_c2_r[16] , \mul_a1/fa1_c2_r[15] , \mul_a1/fa1_c2_r[14] ,
         \mul_a1/fa1_s2_r[33] , \mul_a1/fa1_s2_r[32] , \mul_a1/fa1_s2_r[31] ,
         \mul_a1/fa1_s2_r[30] , \mul_a1/fa1_s2_r[29] , \mul_a1/fa1_s2_r[28] ,
         \mul_a1/fa1_s2_r[27] , \mul_a1/fa1_s2_r[26] , \mul_a1/fa1_s2_r[25] ,
         \mul_a1/fa1_s2_r[24] , \mul_a1/fa1_s2_r[23] , \mul_a1/fa1_s2_r[22] ,
         \mul_a1/fa1_s2_r[21] , \mul_a1/fa1_s2_r[20] , \mul_a1/fa1_s2_r[19] ,
         \mul_a1/fa1_s2_r[18] , \mul_a1/fa1_s2_r[17] , \mul_a1/fa1_s2_r[16] ,
         \mul_a1/fa1_s2_r[15] , \mul_a1/fa1_s2_r[14] , \mul_a1/fa1_s2_r[13] ,
         \mul_a1/fa1_s1_r[33] , \mul_a1/fa1_s1_r[32] , \mul_a1/fa1_s1_r[31] ,
         \mul_a1/fa1_s1_r[30] , \mul_a1/fa1_s1_r[29] , \mul_a1/fa1_s1_r[28] ,
         \mul_a1/fa1_s1_r[27] , \mul_a1/fa1_s1_r[26] , \mul_a1/fa1_s1_r[25] ,
         \mul_a1/fa1_s1_r[24] , \mul_a1/fa1_s1_r[23] , \mul_a1/fa1_s1_r[22] ,
         \mul_a1/fa1_s1_r[21] , \mul_a1/fa1_s1_r[20] , \mul_a1/fa1_s1_r[19] ,
         \mul_a1/fa1_s1_r[18] , \mul_a1/fa1_s1_r[17] , \mul_a1/fa1_s1_r[16] ,
         \mul_a1/fa1_s1_r[15] , \mul_a1/fa1_s1_r[14] , \mul_a1/fa1_s1_r[13] ,
         \mul_a1/fa1_s1_r[12] , \mul_a1/fa1_s1_r[11] , \mul_a1/fa1_s1_r[10] ,
         \mul_a1/fa1_s1_r[9] , \mul_a1/fa1_s1_r[8] , \mul_a1/fa1_c0_r[20] ,
         \mul_a1/fa1_c0_r[19] , \mul_a1/fa1_c0_r[18] , \mul_a1/fa1_c0_r[17] ,
         \mul_a1/fa1_c0_r[16] , \mul_a1/fa1_c0_r[15] , \mul_a1/fa1_c0_r[14] ,
         \mul_a1/fa1_c0_r[13] , \mul_a1/fa1_c0_r[12] , \mul_a1/fa1_c0_r[11] ,
         \mul_a1/fa1_c0_r[10] , \mul_a1/fa1_c0_r[9] , \mul_a1/fa1_c0_r[8] ,
         \mul_a1/fa1_c0_r[7] , \mul_a1/fa1_c0_r[6] , \mul_a1/fa1_c0_r[5] ,
         \mul_a1/fa1_s0_r[33] , \mul_a1/fa1_s0_r[32] , \mul_a1/fa1_s0_r[31] ,
         \mul_a1/fa1_s0_r[30] , \mul_a1/fa1_s0_r[29] , \mul_a1/fa1_s0_r[28] ,
         \mul_a1/fa1_s0_r[27] , \mul_a1/fa1_s0_r[26] , \mul_a1/fa1_s0_r[25] ,
         \mul_a1/fa1_s0_r[24] , \mul_a1/fa1_s0_r[23] , \mul_a1/fa1_s0_r[22] ,
         \mul_a1/fa1_s0_r[21] , \mul_a1/fa1_s0_r[20] , \mul_a1/fa1_s0_r[19] ,
         \mul_a1/fa1_s0_r[18] , \mul_a1/fa1_s0_r[17] , \mul_a1/fa1_s0_r[16] ,
         \mul_a1/fa1_s0_r[15] , \mul_a1/fa1_s0_r[14] , \mul_a1/fa1_s0_r[13] ,
         \mul_a1/fa1_s0_r[12] , \mul_a1/fa1_s0_r[11] , \mul_a1/fa1_s0_r[10] ,
         \mul_a1/fa1_s0_r[9] , \mul_a1/fa1_s0_r[8] , \mul_a1/fa1_s0_r[7] ,
         \mul_a1/fa1_s0_r[6] , \mul_a1/fa1_c2[29] , \mul_a1/fa1_c2[28] ,
         \mul_a1/fa1_c2[27] , \mul_a1/fa1_c2[26] , \mul_a1/fa1_c2[25] ,
         \mul_a1/fa1_c2[24] , \mul_a1/fa1_c2[23] , \mul_a1/fa1_c2[22] ,
         \mul_a1/fa1_c2[21] , \mul_a1/fa1_c2[20] , \mul_a1/fa1_c2[19] ,
         \mul_a1/fa1_c2[18] , \mul_a1/fa1_c2[17] , \mul_a1/fa1_c2[16] ,
         \mul_a1/fa1_c2[15] , \mul_a1/fa1_c2[14] , \mul_a1/fa1_s2[31] ,
         \mul_a1/fa1_s2[30] , \mul_a1/fa1_s2[29] , \mul_a1/fa1_s2[28] ,
         \mul_a1/fa1_s2[27] , \mul_a1/fa1_s2[26] , \mul_a1/fa1_s2[25] ,
         \mul_a1/fa1_s2[24] , \mul_a1/fa1_s2[23] , \mul_a1/fa1_s2[22] ,
         \mul_a1/fa1_s2[21] , \mul_a1/fa1_s2[20] , \mul_a1/fa1_s2[19] ,
         \mul_a1/fa1_s2[18] , \mul_a1/fa1_s2[17] , \mul_a1/fa1_s2[16] ,
         \mul_a1/fa1_s2[15] , \mul_a1/fa1_s2[14] , \mul_a1/fa1_c0[20] ,
         \mul_a1/fa1_c0[19] , \mul_a1/fa1_c0[18] , \mul_a1/fa1_c0[17] ,
         \mul_a1/fa1_c0[16] , \mul_a1/fa1_c0[15] , \mul_a1/fa1_c0[14] ,
         \mul_a1/fa1_c0[13] , \mul_a1/fa1_c0[12] , \mul_a1/fa1_c0[11] ,
         \mul_a1/fa1_c0[10] , \mul_a1/fa1_c0[9] , \mul_a1/fa1_c0[8] ,
         \mul_a1/fa1_c0[7] , \mul_a1/fa1_c0[6] , \mul_a1/fa1_c0[5] ,
         \mul_a1/fa1_s0[27] , \mul_a1/fa1_s0[20] , \mul_a1/fa1_s0[19] ,
         \mul_a1/fa1_s0[18] , \mul_a1/fa1_s0[17] , \mul_a1/fa1_s0[16] ,
         \mul_a1/fa1_s0[15] , \mul_a1/fa1_s0[14] , \mul_a1/fa1_s0[13] ,
         \mul_a1/fa1_s0[12] , \mul_a1/fa1_s0[11] , \mul_a1/fa1_s0[10] ,
         \mul_a1/fa1_s0[9] , \mul_a1/fa1_s0[8] , \mul_a1/fa1_s0[7] ,
         \mul_a1/fa1_s0[6] , \mul_a2/result_sat[15] , \mul_a2/result_sat[14] ,
         \mul_a2/result_sat[13] , \mul_a2/result_sat[12] ,
         \mul_a2/result_sat[11] , \mul_a2/result_sat[10] ,
         \mul_a2/result_sat[9] , \mul_a2/result_sat[8] ,
         \mul_a2/result_sat[7] , \mul_a2/result_sat[6] ,
         \mul_a2/result_sat[5] , \mul_a2/result_sat[4] ,
         \mul_a2/result_sat[3] , \mul_a2/result_sat[2] ,
         \mul_a2/result_sat[1] , \mul_a2/result_sat[0] , \mul_a2/fa1_c2_r[28] ,
         \mul_a2/fa1_c2_r[27] , \mul_a2/fa1_c2_r[26] , \mul_a2/fa1_c2_r[25] ,
         \mul_a2/fa1_c2_r[24] , \mul_a2/fa1_c2_r[23] , \mul_a2/fa1_c2_r[22] ,
         \mul_a2/fa1_c2_r[21] , \mul_a2/fa1_c2_r[20] , \mul_a2/fa1_c2_r[19] ,
         \mul_a2/fa1_c2_r[18] , \mul_a2/fa1_c2_r[17] , \mul_a2/fa1_c2_r[16] ,
         \mul_a2/fa1_c2_r[15] , \mul_a2/fa1_c2_r[14] , \mul_a2/fa1_s2_r[33] ,
         \mul_a2/fa1_s2_r[32] , \mul_a2/fa1_s2_r[31] , \mul_a2/fa1_s2_r[30] ,
         \mul_a2/fa1_s2_r[29] , \mul_a2/fa1_s2_r[28] , \mul_a2/fa1_s2_r[27] ,
         \mul_a2/fa1_s2_r[26] , \mul_a2/fa1_s2_r[25] , \mul_a2/fa1_s2_r[24] ,
         \mul_a2/fa1_s2_r[23] , \mul_a2/fa1_s2_r[22] , \mul_a2/fa1_s2_r[21] ,
         \mul_a2/fa1_s2_r[20] , \mul_a2/fa1_s2_r[19] , \mul_a2/fa1_s2_r[18] ,
         \mul_a2/fa1_s2_r[17] , \mul_a2/fa1_s2_r[16] , \mul_a2/fa1_s2_r[15] ,
         \mul_a2/fa1_s2_r[14] , \mul_a2/fa1_s2_r[13] , \mul_a2/fa1_c1_r[32] ,
         \mul_a2/fa1_c1_r[31] , \mul_a2/fa1_c1_r[30] , \mul_a2/fa1_c1_r[29] ,
         \mul_a2/fa1_c1_r[28] , \mul_a2/fa1_c1_r[27] , \mul_a2/fa1_c1_r[26] ,
         \mul_a2/fa1_c1_r[25] , \mul_a2/fa1_c1_r[24] , \mul_a2/fa1_c1_r[23] ,
         \mul_a2/fa1_c1_r[22] , \mul_a2/fa1_c1_r[21] , \mul_a2/fa1_c1_r[20] ,
         \mul_a2/fa1_c1_r[19] , \mul_a2/fa1_c1_r[18] , \mul_a2/fa1_c1_r[17] ,
         \mul_a2/fa1_c1_r[16] , \mul_a2/fa1_c1_r[15] , \mul_a2/fa1_c1_r[14] ,
         \mul_a2/fa1_c1_r[13] , \mul_a2/fa1_c1_r[12] , \mul_a2/fa1_c1_r[11] ,
         \mul_a2/fa1_c1_r[10] , \mul_a2/fa1_c1_r[9] , \mul_a2/fa1_c1_r[8] ,
         \mul_a2/fa1_s1_r[33] , \mul_a2/fa1_s1_r[32] , \mul_a2/fa1_s1_r[31] ,
         \mul_a2/fa1_s1_r[30] , \mul_a2/fa1_s1_r[29] , \mul_a2/fa1_s1_r[28] ,
         \mul_a2/fa1_s1_r[27] , \mul_a2/fa1_s1_r[26] , \mul_a2/fa1_s1_r[25] ,
         \mul_a2/fa1_s1_r[24] , \mul_a2/fa1_s1_r[23] , \mul_a2/fa1_s1_r[22] ,
         \mul_a2/fa1_s1_r[21] , \mul_a2/fa1_s1_r[20] , \mul_a2/fa1_s1_r[19] ,
         \mul_a2/fa1_s1_r[18] , \mul_a2/fa1_s1_r[17] , \mul_a2/fa1_s1_r[16] ,
         \mul_a2/fa1_s1_r[15] , \mul_a2/fa1_s1_r[14] , \mul_a2/fa1_s1_r[13] ,
         \mul_a2/fa1_s1_r[12] , \mul_a2/fa1_s1_r[11] , \mul_a2/fa1_s1_r[10] ,
         \mul_a2/fa1_s1_r[9] , \mul_a2/fa1_s1_r[8] , \mul_a2/fa1_s1_r[7] ,
         \mul_a2/fa1_s1_r[6] , \mul_a2/fa1_c0_r[32] , \mul_a2/fa1_c0_r[31] ,
         \mul_a2/fa1_c0_r[30] , \mul_a2/fa1_c0_r[29] , \mul_a2/fa1_c0_r[28] ,
         \mul_a2/fa1_c0_r[27] , \mul_a2/fa1_c0_r[26] , \mul_a2/fa1_c0_r[25] ,
         \mul_a2/fa1_c0_r[24] , \mul_a2/fa1_c0_r[23] , \mul_a2/fa1_c0_r[22] ,
         \mul_a2/fa1_c0_r[21] , \mul_a2/fa1_c0_r[20] , \mul_a2/fa1_c0_r[19] ,
         \mul_a2/fa1_c0_r[18] , \mul_a2/fa1_c0_r[17] , \mul_a2/fa1_c0_r[16] ,
         \mul_a2/fa1_c0_r[15] , \mul_a2/fa1_c0_r[14] , \mul_a2/fa1_c0_r[13] ,
         \mul_a2/fa1_c0_r[12] , \mul_a2/fa1_c0_r[11] , \mul_a2/fa1_c0_r[10] ,
         \mul_a2/fa1_c0_r[9] , \mul_a2/fa1_c0_r[8] , \mul_a2/fa1_c0_r[7] ,
         \mul_a2/fa1_c0_r[6] , \mul_a2/fa1_c0_r[5] , \mul_a2/fa1_c0_r[4] ,
         \mul_a2/fa1_c0_r[3] , \mul_a2/fa1_c0_r[2] , \mul_a2/fa1_s0_r[33] ,
         \mul_a2/fa1_s0_r[32] , \mul_a2/fa1_s0_r[31] , \mul_a2/fa1_s0_r[30] ,
         \mul_a2/fa1_s0_r[29] , \mul_a2/fa1_s0_r[28] , \mul_a2/fa1_s0_r[27] ,
         \mul_a2/fa1_s0_r[26] , \mul_a2/fa1_s0_r[25] , \mul_a2/fa1_s0_r[24] ,
         \mul_a2/fa1_s0_r[23] , \mul_a2/fa1_s0_r[22] , \mul_a2/fa1_s0_r[21] ,
         \mul_a2/fa1_s0_r[20] , \mul_a2/fa1_s0_r[19] , \mul_a2/fa1_s0_r[18] ,
         \mul_a2/fa1_s0_r[17] , \mul_a2/fa1_s0_r[16] , \mul_a2/fa1_s0_r[15] ,
         \mul_a2/fa1_s0_r[14] , \mul_a2/fa1_s0_r[13] , \mul_a2/fa1_s0_r[12] ,
         \mul_a2/fa1_s0_r[11] , \mul_a2/fa1_s0_r[10] , \mul_a2/fa1_s0_r[9] ,
         \mul_a2/fa1_s0_r[8] , \mul_a2/fa1_s0_r[7] , \mul_a2/fa1_s0_r[6] ,
         \mul_a2/fa1_s0_r[5] , \mul_a2/fa1_s0_r[4] , \mul_a2/fa1_s0_r[3] ,
         \mul_a2/fa1_c2[28] , \mul_a2/fa1_c2[27] , \mul_a2/fa1_c2[26] ,
         \mul_a2/fa1_c2[25] , \mul_a2/fa1_c2[24] , \mul_a2/fa1_c2[23] ,
         \mul_a2/fa1_c2[22] , \mul_a2/fa1_c2[21] , \mul_a2/fa1_c2[20] ,
         \mul_a2/fa1_c2[19] , \mul_a2/fa1_c2[18] , \mul_a2/fa1_c2[17] ,
         \mul_a2/fa1_c2[16] , \mul_a2/fa1_c2[15] , \mul_a2/fa1_c2[14] ,
         \mul_a2/fa1_s2[31] , \mul_a2/fa1_s2[28] , \mul_a2/fa1_s2[27] ,
         \mul_a2/fa1_s2[26] , \mul_a2/fa1_s2[25] , \mul_a2/fa1_s2[24] ,
         \mul_a2/fa1_s2[23] , \mul_a2/fa1_s2[22] , \mul_a2/fa1_s2[21] ,
         \mul_a2/fa1_s2[20] , \mul_a2/fa1_s2[19] , \mul_a2/fa1_s2[18] ,
         \mul_a2/fa1_s2[17] , \mul_a2/fa1_s2[16] , \mul_a2/fa1_s2[15] ,
         \mul_a2/fa1_s2[14] , \mul_a2/fa1_c1[22] , \mul_a2/fa1_c1[21] ,
         \mul_a2/fa1_c1[20] , \mul_a2/fa1_c1[19] , \mul_a2/fa1_c1[18] ,
         \mul_a2/fa1_c1[17] , \mul_a2/fa1_c1[16] , \mul_a2/fa1_c1[15] ,
         \mul_a2/fa1_c1[14] , \mul_a2/fa1_c1[13] , \mul_a2/fa1_c1[12] ,
         \mul_a2/fa1_c1[11] , \mul_a2/fa1_c1[10] , \mul_a2/fa1_c1[9] ,
         \mul_a2/fa1_c1[8] , \mul_a2/fa1_s1[27] , \mul_a2/fa1_s1[24] ,
         \mul_a2/fa1_s1[23] , \mul_a2/fa1_s1[22] , \mul_a2/fa1_s1[21] ,
         \mul_a2/fa1_s1[20] , \mul_a2/fa1_s1[19] , \mul_a2/fa1_s1[18] ,
         \mul_a2/fa1_s1[17] , \mul_a2/fa1_s1[16] , \mul_a2/fa1_s1[15] ,
         \mul_a2/fa1_s1[14] , \mul_a2/fa1_s1[13] , \mul_a2/fa1_s1[12] ,
         \mul_a2/fa1_s1[11] , \mul_a2/fa1_s1[10] , \mul_a2/fa1_s1[9] ,
         \mul_a2/fa1_s1[8] , \mul_a2/fa1_s1[7] , \mul_a2/fa1_c0[18] ,
         \mul_a2/fa1_c0[17] , \mul_a2/fa1_c0[16] , \mul_a2/fa1_c0[15] ,
         \mul_a2/fa1_c0[14] , \mul_a2/fa1_c0[13] , \mul_a2/fa1_c0[12] ,
         \mul_a2/fa1_c0[11] , \mul_a2/fa1_c0[10] , \mul_a2/fa1_c0[9] ,
         \mul_a2/fa1_c0[8] , \mul_a2/fa1_c0[7] , \mul_a2/fa1_c0[6] ,
         \mul_a2/fa1_c0[5] , \mul_a2/fa1_c0[4] , \mul_a2/fa1_s0[27] ,
         \mul_a2/fa1_s0[20] , \mul_a2/fa1_s0[19] , \mul_a2/fa1_s0[18] ,
         \mul_a2/fa1_s0[17] , \mul_a2/fa1_s0[16] , \mul_a2/fa1_s0[15] ,
         \mul_a2/fa1_s0[14] , \mul_a2/fa1_s0[13] , \mul_a2/fa1_s0[12] ,
         \mul_a2/fa1_s0[11] , \mul_a2/fa1_s0[10] , \mul_a2/fa1_s0[9] ,
         \mul_a2/fa1_s0[8] , \mul_a2/fa1_s0[7] , \mul_a2/fa1_s0[6] ,
         \mul_a2/fa1_s0[5] , \mul_a2/fa1_s0[4] , \mul_a2/fa1_s0[3] ,
         \mul_a2/fa1_s0[1] , \mul_a2/fa1_s0[0] , \C53/DATA4_9 , \C53/DATA4_10 ,
         \C53/DATA4_11 , \C53/DATA4_12 , \C53/DATA4_13 , \C53/DATA4_14 ,
         \C53/DATA4_15 , \C53/DATA4_16 , \C53/DATA4_17 , \C53/DATA4_18 ,
         \C53/DATA4_19 , \C53/DATA4_20 , \C53/DATA4_21 , \C53/DATA4_22 ,
         \C53/DATA4_23 , \C53/DATA4_24 , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988;
  wire   [15:0] x_z1;
  wire   [15:0] x_z2;
  wire   [15:0] y_z1;
  wire   [15:0] y_z2;
  wire   [15:0] x_reg2;
  wire   [15:0] p_b0;
  wire   [15:0] p_b1;
  wire   [15:0] p_b2;
  wire   [15:0] p_a1;
  wire   [15:0] p_a2;

  HS65_GS_DFPRQX4 valid_T1_reg ( .D(n1892), .CP(clk), .RN(rst_n), .Q(valid_T1)
         );
  HS65_GS_DFPRQX4 valid_T2_reg ( .D(valid_T1), .CP(clk), .RN(rst_n), .Q(
        valid_T2) );
  HS65_GS_DFPRQX4 valid_T3_reg ( .D(valid_T2), .CP(clk), .RN(rst_n), .Q(
        valid_T3) );
  HS65_GS_DFPRQX4 valid_out_reg ( .D(valid_T3), .CP(clk), .RN(rst_n), .Q(
        valid_out) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[0]  ( .D(\mul_b0/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[0]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[1]  ( .D(\mul_b0/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[1]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[2]  ( .D(\mul_b0/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[2]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[3]  ( .D(\mul_b0/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[3]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[4]  ( .D(\mul_b0/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[4]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[5]  ( .D(\mul_b0/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[5]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[6]  ( .D(\mul_b0/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[6]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[7]  ( .D(\mul_b0/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[7]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[8]  ( .D(\mul_b0/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[8]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[9]  ( .D(\mul_b0/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[9]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[10]  ( .D(\mul_b0/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[10]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[11]  ( .D(\mul_b0/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[11]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[12]  ( .D(\mul_b0/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[12]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[13]  ( .D(\mul_b0/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[13]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[14]  ( .D(\mul_b0/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[14]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[15]  ( .D(\mul_b0/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[15]) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[12]  ( .D(x_z1[0]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[13]  ( .D(x_z1[1]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[14]  ( .D(x_z1[2]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[15]  ( .D(x_z1[3]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[16]  ( .D(x_z1[4]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[17]  ( .D(x_z1[5]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[18]  ( .D(x_z1[6]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[19]  ( .D(x_z1[7]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[20]  ( .D(x_z1[8]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[21]  ( .D(x_z1[9]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[22]  ( .D(x_z1[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[23]  ( .D(x_z1[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[24]  ( .D(x_z1[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[25]  ( .D(x_z1[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[26]  ( .D(x_z1[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[27]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[28]  ( .D(n1891), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[29]  ( .D(n1891), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[30]  ( .D(n1891), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[31]  ( .D(n1891), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[32]  ( .D(n1891), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[33]  ( .D(n1891), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[8]  ( .D(x_z1[0]), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[9]  ( .D(x_z1[1]), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[10]  ( .D(x_z1[2]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[11]  ( .D(x_z1[3]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[12]  ( .D(x_z1[4]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[13]  ( .D(x_z1[5]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[14]  ( .D(x_z1[6]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[15]  ( .D(x_z1[7]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[16]  ( .D(x_z1[8]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[17]  ( .D(x_z1[9]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[18]  ( .D(x_z1[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[19]  ( .D(x_z1[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[20]  ( .D(x_z1[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[21]  ( .D(x_z1[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[22]  ( .D(x_z1[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[23]  ( .D(n1891), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[24]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[25]  ( .D(n1891), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[26]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[27]  ( .D(n1891), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[28]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[29]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[30]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[31]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[32]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[33]  ( .D(n1891), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[5]  ( .D(\mul_b0/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[6]  ( .D(\mul_b0/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[7]  ( .D(\mul_b0/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[8]  ( .D(\mul_b0/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[9]  ( .D(\mul_b0/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[10]  ( .D(\mul_b0/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[11]  ( .D(\mul_b0/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[12]  ( .D(\mul_b0/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[13]  ( .D(\mul_b0/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[14]  ( .D(\mul_b0/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[15]  ( .D(\mul_b0/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[16]  ( .D(\mul_b0/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[17]  ( .D(\mul_b0/fa1_c0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[18]  ( .D(\mul_b0/fa1_c0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[19]  ( .D(\mul_b0/fa1_c0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[20]  ( .D(\mul_b0/fa1_c0[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[6]  ( .D(\mul_b0/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[7]  ( .D(\mul_b0/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[8]  ( .D(\mul_b0/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[9]  ( .D(\mul_b0/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[10]  ( .D(\mul_b0/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[11]  ( .D(\mul_b0/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[12]  ( .D(\mul_b0/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[13]  ( .D(\mul_b0/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[14]  ( .D(\mul_b0/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[15]  ( .D(\mul_b0/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[16]  ( .D(\mul_b0/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[17]  ( .D(\mul_b0/fa1_s0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[18]  ( .D(\mul_b0/fa1_s0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[19]  ( .D(\mul_b0/fa1_s0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[20]  ( .D(\mul_b0/fa1_s0[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[21]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[22]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[23]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[24]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[25]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[26]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[27]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[28]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[29]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[30]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[31]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[32]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[33]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[0]  ( .D(\mul_b1/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[0]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[1]  ( .D(\mul_b1/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[1]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[2]  ( .D(\mul_b1/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[2]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[3]  ( .D(\mul_b1/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[3]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[4]  ( .D(\mul_b1/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[4]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[5]  ( .D(\mul_b1/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[5]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[6]  ( .D(\mul_b1/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[6]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[7]  ( .D(\mul_b1/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[7]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[8]  ( .D(\mul_b1/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[8]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[9]  ( .D(\mul_b1/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[9]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[10]  ( .D(\mul_b1/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[10]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[11]  ( .D(\mul_b1/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[11]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[12]  ( .D(\mul_b1/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[12]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[13]  ( .D(\mul_b1/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[13]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[14]  ( .D(\mul_b1/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[14]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[15]  ( .D(\mul_b1/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[15]) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[13]  ( .D(x_z2[0]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[14]  ( .D(\mul_b1/fa1_s2[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[15]  ( .D(\mul_b1/fa1_s2[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[16]  ( .D(\mul_b1/fa1_s2[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[17]  ( .D(\mul_b1/fa1_s2[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[18]  ( .D(\mul_b1/fa1_s2[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[19]  ( .D(\mul_b1/fa1_s2[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[20]  ( .D(\mul_b1/fa1_s2[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[21]  ( .D(\mul_b1/fa1_s2[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[22]  ( .D(\mul_b1/fa1_s2[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[23]  ( .D(\mul_b1/fa1_s2[23] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[24]  ( .D(\mul_b1/fa1_s2[24] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[25]  ( .D(\mul_b1/fa1_s2[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[26]  ( .D(\mul_b1/fa1_s2[26] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[27]  ( .D(\mul_b1/fa1_s2[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[28]  ( .D(\mul_b1/fa1_s2[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[29]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[30]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[31]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[32]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[33]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[9]  ( .D(x_z2[0]), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[10]  ( .D(x_z2[1]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[11]  ( .D(x_z2[2]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[12]  ( .D(x_z2[3]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[13]  ( .D(x_z2[4]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[14]  ( .D(x_z2[5]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[15]  ( .D(x_z2[6]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[16]  ( .D(x_z2[7]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[17]  ( .D(x_z2[8]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[18]  ( .D(x_z2[9]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[19]  ( .D(x_z2[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[20]  ( .D(x_z2[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[21]  ( .D(x_z2[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[22]  ( .D(x_z2[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[23]  ( .D(x_z2[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[24]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[25]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[26]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[27]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[28]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[29]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[30]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[31]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[32]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[33]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[4]  ( .D(\mul_b1/fa1_c0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[5]  ( .D(\mul_b1/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[6]  ( .D(\mul_b1/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[7]  ( .D(\mul_b1/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[8]  ( .D(\mul_b1/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[9]  ( .D(\mul_b1/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[10]  ( .D(\mul_b1/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[11]  ( .D(\mul_b1/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[12]  ( .D(\mul_b1/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[13]  ( .D(\mul_b1/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[14]  ( .D(\mul_b1/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[15]  ( .D(\mul_b1/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[16]  ( .D(\mul_b1/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[17]  ( .D(\mul_b1/fa1_c0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[18]  ( .D(\mul_b1/fa1_c0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[19]  ( .D(\mul_b1/fa1_c0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[5]  ( .D(\mul_b1/fa1_s0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[6]  ( .D(\mul_b1/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[7]  ( .D(\mul_b1/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[8]  ( .D(\mul_b1/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[9]  ( .D(\mul_b1/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[10]  ( .D(\mul_b1/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[11]  ( .D(\mul_b1/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[12]  ( .D(\mul_b1/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[13]  ( .D(\mul_b1/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[14]  ( .D(\mul_b1/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[15]  ( .D(\mul_b1/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[16]  ( .D(\mul_b1/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[17]  ( .D(\mul_b1/fa1_s0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[18]  ( .D(\mul_b1/fa1_s0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[19]  ( .D(\mul_b1/fa1_s0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[20]  ( .D(\mul_b1/fa1_s0[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[21]  ( .D(\mul_b1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[22]  ( .D(\mul_b1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[23]  ( .D(\mul_b1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[24]  ( .D(\mul_b1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[25]  ( .D(\mul_b1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[26]  ( .D(\mul_b1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[27]  ( .D(\mul_b1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[28]  ( .D(\mul_b1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[29]  ( .D(\mul_b1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[30]  ( .D(\mul_b1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[31]  ( .D(\mul_b1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[32]  ( .D(\mul_b1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[33]  ( .D(\mul_b1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[14]  ( .D(\mul_b1/fa1_c2[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[15]  ( .D(\mul_b1/fa1_c2[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[16]  ( .D(\mul_b1/fa1_c2[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[17]  ( .D(\mul_b1/fa1_c2[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[18]  ( .D(\mul_b1/fa1_c2[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[19]  ( .D(\mul_b1/fa1_c2[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[20]  ( .D(\mul_b1/fa1_c2[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[21]  ( .D(\mul_b1/fa1_c2[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[22]  ( .D(\mul_b1/fa1_c2[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[23]  ( .D(\mul_b1/fa1_c2[23] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[24]  ( .D(\mul_b1/fa1_c2[24] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[25]  ( .D(\mul_b1/fa1_c2[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[26]  ( .D(\mul_b1/fa1_c2[26] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[27]  ( .D(\mul_b1/fa1_c2[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[28]  ( .D(\mul_b1/fa1_c2[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[0]  ( .D(\mul_b2/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[0]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[1]  ( .D(\mul_b2/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[1]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[2]  ( .D(\mul_b2/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[2]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[3]  ( .D(\mul_b2/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[3]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[4]  ( .D(\mul_b2/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[4]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[5]  ( .D(\mul_b2/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[5]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[6]  ( .D(\mul_b2/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[6]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[7]  ( .D(\mul_b2/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[7]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[8]  ( .D(\mul_b2/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[8]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[9]  ( .D(\mul_b2/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[9]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[10]  ( .D(\mul_b2/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[10]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[11]  ( .D(\mul_b2/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[11]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[12]  ( .D(\mul_b2/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[12]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[13]  ( .D(\mul_b2/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[13]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[14]  ( .D(\mul_b2/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[14]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[15]  ( .D(\mul_b2/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[15]) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[12]  ( .D(x_reg2[0]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[13]  ( .D(x_reg2[1]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[14]  ( .D(x_reg2[2]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[15]  ( .D(x_reg2[3]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[16]  ( .D(x_reg2[4]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[17]  ( .D(x_reg2[5]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[18]  ( .D(x_reg2[6]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[19]  ( .D(x_reg2[7]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[20]  ( .D(x_reg2[8]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[21]  ( .D(x_reg2[9]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[22]  ( .D(x_reg2[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[23]  ( .D(x_reg2[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[24]  ( .D(x_reg2[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[25]  ( .D(x_reg2[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[26]  ( .D(x_reg2[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[27]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[28]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[29]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[30]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[31]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[32]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[33]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[8]  ( .D(x_reg2[0]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[9]  ( .D(x_reg2[1]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[10]  ( .D(x_reg2[2]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[11]  ( .D(x_reg2[3]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[12]  ( .D(x_reg2[4]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[13]  ( .D(x_reg2[5]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[14]  ( .D(x_reg2[6]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[15]  ( .D(x_reg2[7]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[16]  ( .D(x_reg2[8]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[17]  ( .D(x_reg2[9]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[18]  ( .D(x_reg2[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[19]  ( .D(x_reg2[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[20]  ( .D(x_reg2[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[21]  ( .D(x_reg2[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[22]  ( .D(x_reg2[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[23]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[24]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[25]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[26]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[27]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[28]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[29]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[30]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[31]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[32]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[33]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[2]  ( .D(\mul_b2/fa1_c0[2] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[2] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[3]  ( .D(\mul_b2/fa1_c0[3] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[3] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[4]  ( .D(\mul_b2/fa1_c0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[5]  ( .D(\mul_b2/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[6]  ( .D(\mul_b2/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[7]  ( .D(\mul_b2/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[8]  ( .D(\mul_b2/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[9]  ( .D(\mul_b2/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[10]  ( .D(\mul_b2/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[11]  ( .D(\mul_b2/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[12]  ( .D(\mul_b2/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[13]  ( .D(\mul_b2/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[14]  ( .D(\mul_b2/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[15]  ( .D(\mul_b2/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[16]  ( .D(\mul_b2/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[17]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[18]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[19]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[20]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[21]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[22]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[23]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[24]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[25]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[26]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[27]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[28]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[29]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[30]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[31]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[32]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[3]  ( .D(\mul_b2/fa1_s0[3] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[3] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[4]  ( .D(\mul_b2/fa1_s0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[5]  ( .D(\mul_b2/fa1_s0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[6]  ( .D(\mul_b2/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[7]  ( .D(\mul_b2/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[8]  ( .D(\mul_b2/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[9]  ( .D(\mul_b2/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[10]  ( .D(\mul_b2/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[11]  ( .D(\mul_b2/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[12]  ( .D(\mul_b2/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[13]  ( .D(\mul_b2/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[14]  ( .D(\mul_b2/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[15]  ( .D(\mul_b2/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[16]  ( .D(\mul_b2/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[17]  ( .D(x_reg2[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[18]  ( .D(x_reg2[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[19]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[20]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[21]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[22]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[23]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[24]  ( .D(n1890), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[25]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[26]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[27]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[28]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[29]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[30]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[31]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[32]  ( .D(n1889), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[33]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[0]  ( .D(\mul_a1/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[0]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[1]  ( .D(\mul_a1/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[1]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[2]  ( .D(\mul_a1/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[2]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[3]  ( .D(\mul_a1/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[3]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[4]  ( .D(\mul_a1/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[4]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[5]  ( .D(\mul_a1/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[5]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[6]  ( .D(\mul_a1/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[6]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[7]  ( .D(\mul_a1/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[7]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[8]  ( .D(\mul_a1/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[8]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[9]  ( .D(\mul_a1/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[9]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[10]  ( .D(\mul_a1/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[10]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[11]  ( .D(\mul_a1/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[11]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[12]  ( .D(\mul_a1/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[12]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[13]  ( .D(\mul_a1/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[13]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[14]  ( .D(\mul_a1/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[14]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[15]  ( .D(\mul_a1/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[15]) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[13]  ( .D(y_z1[0]), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[14]  ( .D(\mul_a1/fa1_s2[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[15]  ( .D(\mul_a1/fa1_s2[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[16]  ( .D(\mul_a1/fa1_s2[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[17]  ( .D(\mul_a1/fa1_s2[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[18]  ( .D(\mul_a1/fa1_s2[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[19]  ( .D(\mul_a1/fa1_s2[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[20]  ( .D(\mul_a1/fa1_s2[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[21]  ( .D(\mul_a1/fa1_s2[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[22]  ( .D(\mul_a1/fa1_s2[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[23]  ( .D(\mul_a1/fa1_s2[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[24]  ( .D(\mul_a1/fa1_s2[24] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[25]  ( .D(\mul_a1/fa1_s2[25] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[26]  ( .D(\mul_a1/fa1_s2[26] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[27]  ( .D(\mul_a1/fa1_s2[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[28]  ( .D(\mul_a1/fa1_s2[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[29]  ( .D(\mul_a1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[30]  ( .D(\mul_a1/fa1_s2[30] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[31]  ( .D(\mul_a1/fa1_s2[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[32]  ( .D(\mul_a1/fa1_s2[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[33]  ( .D(\mul_a1/fa1_s2[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[8]  ( .D(y_z1[0]), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[9]  ( .D(\C53/DATA4_9 ), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[10]  ( .D(\C53/DATA4_10 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[11]  ( .D(\C53/DATA4_11 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[12]  ( .D(\C53/DATA4_12 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[13]  ( .D(\C53/DATA4_13 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[14]  ( .D(\C53/DATA4_14 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[15]  ( .D(\C53/DATA4_15 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[16]  ( .D(\C53/DATA4_16 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[17]  ( .D(\C53/DATA4_17 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[18]  ( .D(\C53/DATA4_18 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[19]  ( .D(\C53/DATA4_19 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[20]  ( .D(\C53/DATA4_20 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[21]  ( .D(\C53/DATA4_21 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[22]  ( .D(\C53/DATA4_22 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[23]  ( .D(\C53/DATA4_23 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[24]  ( .D(\C53/DATA4_24 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[25]  ( .D(n1886), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[26]  ( .D(n1886), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[27]  ( .D(n1886), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[28]  ( .D(n1886), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[29]  ( .D(n1886), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[30]  ( .D(n1886), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[31]  ( .D(n1886), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[32]  ( .D(n1886), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[33]  ( .D(n1886), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[5]  ( .D(\mul_a1/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[6]  ( .D(\mul_a1/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[7]  ( .D(\mul_a1/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[8]  ( .D(\mul_a1/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[9]  ( .D(\mul_a1/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[10]  ( .D(\mul_a1/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[11]  ( .D(\mul_a1/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[12]  ( .D(\mul_a1/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[13]  ( .D(\mul_a1/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[14]  ( .D(\mul_a1/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[15]  ( .D(\mul_a1/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[16]  ( .D(\mul_a1/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[17]  ( .D(\mul_a1/fa1_c0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[18]  ( .D(\mul_a1/fa1_c0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[19]  ( .D(\mul_a1/fa1_c0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[20]  ( .D(\mul_a1/fa1_c0[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[6]  ( .D(\mul_a1/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[7]  ( .D(\mul_a1/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[8]  ( .D(\mul_a1/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[9]  ( .D(\mul_a1/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[10]  ( .D(\mul_a1/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[11]  ( .D(\mul_a1/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[12]  ( .D(\mul_a1/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[13]  ( .D(\mul_a1/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[14]  ( .D(\mul_a1/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[15]  ( .D(\mul_a1/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[16]  ( .D(\mul_a1/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[17]  ( .D(\mul_a1/fa1_s0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[18]  ( .D(\mul_a1/fa1_s0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[19]  ( .D(\mul_a1/fa1_s0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[20]  ( .D(\mul_a1/fa1_s0[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[21]  ( .D(\mul_a1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[22]  ( .D(\mul_a1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[23]  ( .D(\mul_a1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[24]  ( .D(\mul_a1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[25]  ( .D(\mul_a1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[26]  ( .D(\mul_a1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[27]  ( .D(\mul_a1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[28]  ( .D(\mul_a1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[29]  ( .D(\mul_a1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[30]  ( .D(\mul_a1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[31]  ( .D(\mul_a1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[32]  ( .D(\mul_a1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[33]  ( .D(\mul_a1/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[14]  ( .D(\mul_a1/fa1_c2[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[15]  ( .D(\mul_a1/fa1_c2[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[16]  ( .D(\mul_a1/fa1_c2[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[17]  ( .D(\mul_a1/fa1_c2[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[18]  ( .D(\mul_a1/fa1_c2[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[19]  ( .D(\mul_a1/fa1_c2[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[20]  ( .D(\mul_a1/fa1_c2[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[21]  ( .D(\mul_a1/fa1_c2[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[22]  ( .D(\mul_a1/fa1_c2[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[23]  ( .D(\mul_a1/fa1_c2[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[24]  ( .D(\mul_a1/fa1_c2[24] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[25]  ( .D(\mul_a1/fa1_c2[25] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[26]  ( .D(\mul_a1/fa1_c2[26] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[27]  ( .D(\mul_a1/fa1_c2[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[28]  ( .D(\mul_a1/fa1_c2[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[29]  ( .D(\mul_a1/fa1_c2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[0]  ( .D(\mul_a2/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[0]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[1]  ( .D(\mul_a2/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[1]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[2]  ( .D(\mul_a2/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[2]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[3]  ( .D(\mul_a2/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[3]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[4]  ( .D(\mul_a2/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[4]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[5]  ( .D(\mul_a2/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[5]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[6]  ( .D(\mul_a2/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[6]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[7]  ( .D(\mul_a2/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[7]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[8]  ( .D(\mul_a2/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[8]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[9]  ( .D(\mul_a2/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[9]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[10]  ( .D(\mul_a2/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[10]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[11]  ( .D(\mul_a2/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[11]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[12]  ( .D(\mul_a2/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[12]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[13]  ( .D(\mul_a2/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[13]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[14]  ( .D(\mul_a2/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[14]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[15]  ( .D(\mul_a2/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[15]) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[13]  ( .D(\mul_a2/fa1_s0[0] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[14]  ( .D(\mul_a2/fa1_s2[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[15]  ( .D(\mul_a2/fa1_s2[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[16]  ( .D(\mul_a2/fa1_s2[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[17]  ( .D(\mul_a2/fa1_s2[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[18]  ( .D(\mul_a2/fa1_s2[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[19]  ( .D(\mul_a2/fa1_s2[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[20]  ( .D(\mul_a2/fa1_s2[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[21]  ( .D(\mul_a2/fa1_s2[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[22]  ( .D(\mul_a2/fa1_s2[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[23]  ( .D(\mul_a2/fa1_s2[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[24]  ( .D(\mul_a2/fa1_s2[24] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[25]  ( .D(\mul_a2/fa1_s2[25] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[26]  ( .D(\mul_a2/fa1_s2[26] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[27]  ( .D(\mul_a2/fa1_s2[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[28]  ( .D(\mul_a2/fa1_s2[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[29]  ( .D(\mul_a2/fa1_s2[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[30]  ( .D(\mul_a2/fa1_s2[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[31]  ( .D(\mul_a2/fa1_s2[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[32]  ( .D(\mul_a2/fa1_s2[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[33]  ( .D(\mul_a2/fa1_s2[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[8]  ( .D(\mul_a2/fa1_c1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[9]  ( .D(\mul_a2/fa1_c1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[10]  ( .D(\mul_a2/fa1_c1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[11]  ( .D(\mul_a2/fa1_c1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[12]  ( .D(\mul_a2/fa1_c1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[13]  ( .D(\mul_a2/fa1_c1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[14]  ( .D(\mul_a2/fa1_c1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[15]  ( .D(\mul_a2/fa1_c1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[16]  ( .D(\mul_a2/fa1_c1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[17]  ( .D(\mul_a2/fa1_c1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[18]  ( .D(\mul_a2/fa1_c1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[19]  ( .D(\mul_a2/fa1_c1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[20]  ( .D(\mul_a2/fa1_c1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[21]  ( .D(\mul_a2/fa1_c1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[22]  ( .D(\mul_a2/fa1_c1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[23]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[24]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[25]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[26]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[27]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[28]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[29]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[30]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[31]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[32]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[6]  ( .D(\mul_a2/fa1_s0[0] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[6] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[7]  ( .D(\mul_a2/fa1_s1[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[8]  ( .D(\mul_a2/fa1_s1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[9]  ( .D(\mul_a2/fa1_s1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[10]  ( .D(\mul_a2/fa1_s1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[11]  ( .D(\mul_a2/fa1_s1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[12]  ( .D(\mul_a2/fa1_s1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[13]  ( .D(\mul_a2/fa1_s1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[14]  ( .D(\mul_a2/fa1_s1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[15]  ( .D(\mul_a2/fa1_s1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[16]  ( .D(\mul_a2/fa1_s1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[17]  ( .D(\mul_a2/fa1_s1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[18]  ( .D(\mul_a2/fa1_s1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[19]  ( .D(\mul_a2/fa1_s1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[20]  ( .D(\mul_a2/fa1_s1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[21]  ( .D(\mul_a2/fa1_s1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[22]  ( .D(\mul_a2/fa1_s1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[23]  ( .D(\mul_a2/fa1_s1[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[24]  ( .D(\mul_a2/fa1_s1[24] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[25]  ( .D(\mul_a2/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[26]  ( .D(\mul_a2/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[27]  ( .D(\mul_a2/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[28]  ( .D(\mul_a2/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[29]  ( .D(\mul_a2/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[30]  ( .D(\mul_a2/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[31]  ( .D(\mul_a2/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[32]  ( .D(\mul_a2/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[33]  ( .D(\mul_a2/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[2]  ( .D(n1885), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c0_r[2] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[3]  ( .D(n1887), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c0_r[3] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[4]  ( .D(\mul_a2/fa1_c0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[5]  ( .D(\mul_a2/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[6]  ( .D(\mul_a2/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[7]  ( .D(\mul_a2/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[8]  ( .D(\mul_a2/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[9]  ( .D(\mul_a2/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[10]  ( .D(\mul_a2/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[11]  ( .D(\mul_a2/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[12]  ( .D(\mul_a2/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[13]  ( .D(\mul_a2/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[14]  ( .D(\mul_a2/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[15]  ( .D(\mul_a2/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[16]  ( .D(\mul_a2/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[17]  ( .D(\mul_a2/fa1_c0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[18]  ( .D(\mul_a2/fa1_c0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[19]  ( .D(n1888), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[20]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[21]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[22]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[23]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[24]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[25]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[26]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[27]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[28]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[29]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[30]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[31]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[32]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[3]  ( .D(\mul_a2/fa1_s0[3] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[3] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[4]  ( .D(\mul_a2/fa1_s0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[5]  ( .D(\mul_a2/fa1_s0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[6]  ( .D(\mul_a2/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[7]  ( .D(\mul_a2/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[8]  ( .D(\mul_a2/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[9]  ( .D(\mul_a2/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[10]  ( .D(\mul_a2/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[11]  ( .D(\mul_a2/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[12]  ( .D(\mul_a2/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[13]  ( .D(\mul_a2/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[14]  ( .D(\mul_a2/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[15]  ( .D(\mul_a2/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[16]  ( .D(\mul_a2/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[17]  ( .D(\mul_a2/fa1_s0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[18]  ( .D(\mul_a2/fa1_s0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[19]  ( .D(\mul_a2/fa1_s0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[20]  ( .D(\mul_a2/fa1_s0[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[21]  ( .D(\mul_a2/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[22]  ( .D(\mul_a2/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[23]  ( .D(\mul_a2/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[24]  ( .D(\mul_a2/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[25]  ( .D(\mul_a2/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[26]  ( .D(\mul_a2/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[27]  ( .D(\mul_a2/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[28]  ( .D(\mul_a2/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[29]  ( .D(\mul_a2/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[30]  ( .D(\mul_a2/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[31]  ( .D(\mul_a2/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[32]  ( .D(\mul_a2/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[33]  ( .D(\mul_a2/fa1_s0[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[14]  ( .D(\mul_a2/fa1_c2[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[15]  ( .D(\mul_a2/fa1_c2[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[16]  ( .D(\mul_a2/fa1_c2[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[17]  ( .D(\mul_a2/fa1_c2[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[18]  ( .D(\mul_a2/fa1_c2[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[19]  ( .D(\mul_a2/fa1_c2[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[20]  ( .D(\mul_a2/fa1_c2[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[21]  ( .D(\mul_a2/fa1_c2[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[22]  ( .D(\mul_a2/fa1_c2[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[23]  ( .D(\mul_a2/fa1_c2[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[24]  ( .D(\mul_a2/fa1_c2[24] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[25]  ( .D(\mul_a2/fa1_c2[25] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[26]  ( .D(\mul_a2/fa1_c2[26] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[27]  ( .D(\mul_a2/fa1_c2[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[28]  ( .D(\mul_a2/fa1_c2[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[28] ) );
  HS65_GS_DFPRQX4 \x_z1_reg[15]  ( .D(n1893), .CP(clk), .RN(rst_n), .Q(
        x_z1[15]) );
  HS65_GS_DFPRQX4 \x_z1_reg[14]  ( .D(n1894), .CP(clk), .RN(rst_n), .Q(
        x_z1[14]) );
  HS65_GS_DFPRQX4 \x_z1_reg[13]  ( .D(n1895), .CP(clk), .RN(rst_n), .Q(
        x_z1[13]) );
  HS65_GS_DFPRQX4 \x_z1_reg[12]  ( .D(n1896), .CP(clk), .RN(rst_n), .Q(
        x_z1[12]) );
  HS65_GS_DFPRQX4 \x_z1_reg[11]  ( .D(n1897), .CP(clk), .RN(rst_n), .Q(
        x_z1[11]) );
  HS65_GS_DFPRQX4 \x_z1_reg[10]  ( .D(n1898), .CP(clk), .RN(rst_n), .Q(
        x_z1[10]) );
  HS65_GS_DFPRQX4 \x_z1_reg[9]  ( .D(n1899), .CP(clk), .RN(rst_n), .Q(x_z1[9])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[8]  ( .D(n1900), .CP(clk), .RN(rst_n), .Q(x_z1[8])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[7]  ( .D(n1901), .CP(clk), .RN(rst_n), .Q(x_z1[7])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[6]  ( .D(n1902), .CP(clk), .RN(rst_n), .Q(x_z1[6])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[5]  ( .D(n1903), .CP(clk), .RN(rst_n), .Q(x_z1[5])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[4]  ( .D(n1904), .CP(clk), .RN(rst_n), .Q(x_z1[4])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[3]  ( .D(n1905), .CP(clk), .RN(rst_n), .Q(x_z1[3])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[2]  ( .D(n1906), .CP(clk), .RN(rst_n), .Q(x_z1[2])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[1]  ( .D(n1907), .CP(clk), .RN(rst_n), .Q(x_z1[1])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[0]  ( .D(n1908), .CP(clk), .RN(rst_n), .Q(x_z1[0])
         );
  HS65_GS_DFPRQX4 \x_z2_reg[15]  ( .D(n1909), .CP(clk), .RN(rst_n), .Q(
        x_z2[15]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[15]  ( .D(n1910), .CP(clk), .RN(rst_n), .Q(
        x_reg2[15]) );
  HS65_GS_DFPRQX4 \x_z2_reg[14]  ( .D(n1911), .CP(clk), .RN(rst_n), .Q(
        x_z2[14]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[14]  ( .D(n1912), .CP(clk), .RN(rst_n), .Q(
        x_reg2[14]) );
  HS65_GS_DFPRQX4 \x_z2_reg[13]  ( .D(n1913), .CP(clk), .RN(rst_n), .Q(
        x_z2[13]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[13]  ( .D(n1914), .CP(clk), .RN(rst_n), .Q(
        x_reg2[13]) );
  HS65_GS_DFPRQX4 \x_z2_reg[12]  ( .D(n1915), .CP(clk), .RN(rst_n), .Q(
        x_z2[12]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[12]  ( .D(n1916), .CP(clk), .RN(rst_n), .Q(
        x_reg2[12]) );
  HS65_GS_DFPRQX4 \x_z2_reg[11]  ( .D(n1917), .CP(clk), .RN(rst_n), .Q(
        x_z2[11]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[11]  ( .D(n1918), .CP(clk), .RN(rst_n), .Q(
        x_reg2[11]) );
  HS65_GS_DFPRQX4 \x_z2_reg[10]  ( .D(n1919), .CP(clk), .RN(rst_n), .Q(
        x_z2[10]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[10]  ( .D(n1920), .CP(clk), .RN(rst_n), .Q(
        x_reg2[10]) );
  HS65_GS_DFPRQX4 \x_z2_reg[9]  ( .D(n1921), .CP(clk), .RN(rst_n), .Q(x_z2[9])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[9]  ( .D(n1922), .CP(clk), .RN(rst_n), .Q(
        x_reg2[9]) );
  HS65_GS_DFPRQX4 \x_z2_reg[8]  ( .D(n1923), .CP(clk), .RN(rst_n), .Q(x_z2[8])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[8]  ( .D(n1924), .CP(clk), .RN(rst_n), .Q(
        x_reg2[8]) );
  HS65_GS_DFPRQX4 \x_z2_reg[7]  ( .D(n1925), .CP(clk), .RN(rst_n), .Q(x_z2[7])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[7]  ( .D(n1926), .CP(clk), .RN(rst_n), .Q(
        x_reg2[7]) );
  HS65_GS_DFPRQX4 \x_z2_reg[6]  ( .D(n1927), .CP(clk), .RN(rst_n), .Q(x_z2[6])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[6]  ( .D(n1928), .CP(clk), .RN(rst_n), .Q(
        x_reg2[6]) );
  HS65_GS_DFPRQX4 \x_z2_reg[5]  ( .D(n1929), .CP(clk), .RN(rst_n), .Q(x_z2[5])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[5]  ( .D(n1930), .CP(clk), .RN(rst_n), .Q(
        x_reg2[5]) );
  HS65_GS_DFPRQX4 \x_z2_reg[4]  ( .D(n1931), .CP(clk), .RN(rst_n), .Q(x_z2[4])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[4]  ( .D(n1932), .CP(clk), .RN(rst_n), .Q(
        x_reg2[4]) );
  HS65_GS_DFPRQX4 \x_z2_reg[3]  ( .D(n1933), .CP(clk), .RN(rst_n), .Q(x_z2[3])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[3]  ( .D(n1934), .CP(clk), .RN(rst_n), .Q(
        x_reg2[3]) );
  HS65_GS_DFPRQX4 \x_z2_reg[2]  ( .D(n1935), .CP(clk), .RN(rst_n), .Q(x_z2[2])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[2]  ( .D(n1936), .CP(clk), .RN(rst_n), .Q(
        x_reg2[2]) );
  HS65_GS_DFPRQX4 \x_z2_reg[1]  ( .D(n1937), .CP(clk), .RN(rst_n), .Q(x_z2[1])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[1]  ( .D(n1938), .CP(clk), .RN(rst_n), .Q(
        x_reg2[1]) );
  HS65_GS_DFPRQX4 \x_z2_reg[0]  ( .D(n1939), .CP(clk), .RN(rst_n), .Q(x_z2[0])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[0]  ( .D(n1940), .CP(clk), .RN(rst_n), .Q(
        x_reg2[0]) );
  HS65_GS_DFPRQX4 \data_out_reg[15]  ( .D(n1941), .CP(clk), .RN(rst_n), .Q(
        data_out[15]) );
  HS65_GS_DFPRQX4 \y_z1_reg[15]  ( .D(n1942), .CP(clk), .RN(rst_n), .Q(
        y_z1[15]) );
  HS65_GS_DFPRQX4 \y_z2_reg[15]  ( .D(n1943), .CP(clk), .RN(rst_n), .Q(
        y_z2[15]) );
  HS65_GS_DFPRQX4 \data_out_reg[14]  ( .D(n1944), .CP(clk), .RN(rst_n), .Q(
        data_out[14]) );
  HS65_GS_DFPRQX4 \y_z1_reg[14]  ( .D(n1945), .CP(clk), .RN(rst_n), .Q(
        y_z1[14]) );
  HS65_GS_DFPRQX4 \y_z2_reg[14]  ( .D(n1946), .CP(clk), .RN(rst_n), .Q(
        y_z2[14]) );
  HS65_GS_DFPRQX4 \data_out_reg[13]  ( .D(n1947), .CP(clk), .RN(rst_n), .Q(
        data_out[13]) );
  HS65_GS_DFPRQX4 \y_z1_reg[13]  ( .D(n1948), .CP(clk), .RN(rst_n), .Q(
        y_z1[13]) );
  HS65_GS_DFPRQX4 \y_z2_reg[13]  ( .D(n1949), .CP(clk), .RN(rst_n), .Q(
        y_z2[13]) );
  HS65_GS_DFPRQX4 \data_out_reg[12]  ( .D(n1950), .CP(clk), .RN(rst_n), .Q(
        data_out[12]) );
  HS65_GS_DFPRQX4 \y_z1_reg[12]  ( .D(n1951), .CP(clk), .RN(rst_n), .Q(
        y_z1[12]) );
  HS65_GS_DFPRQX4 \y_z2_reg[12]  ( .D(n1952), .CP(clk), .RN(rst_n), .Q(
        y_z2[12]) );
  HS65_GS_DFPRQX4 \data_out_reg[11]  ( .D(n1953), .CP(clk), .RN(rst_n), .Q(
        data_out[11]) );
  HS65_GS_DFPRQX4 \y_z1_reg[11]  ( .D(n1954), .CP(clk), .RN(rst_n), .Q(
        y_z1[11]) );
  HS65_GS_DFPRQX4 \y_z2_reg[11]  ( .D(n1955), .CP(clk), .RN(rst_n), .Q(
        y_z2[11]) );
  HS65_GS_DFPRQX4 \data_out_reg[10]  ( .D(n1956), .CP(clk), .RN(rst_n), .Q(
        data_out[10]) );
  HS65_GS_DFPRQX4 \y_z1_reg[10]  ( .D(n1957), .CP(clk), .RN(rst_n), .Q(
        y_z1[10]) );
  HS65_GS_DFPRQX4 \y_z2_reg[10]  ( .D(n1958), .CP(clk), .RN(rst_n), .Q(
        y_z2[10]) );
  HS65_GS_DFPRQX4 \data_out_reg[9]  ( .D(n1959), .CP(clk), .RN(rst_n), .Q(
        data_out[9]) );
  HS65_GS_DFPRQX4 \y_z1_reg[9]  ( .D(n1960), .CP(clk), .RN(rst_n), .Q(y_z1[9])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[9]  ( .D(n1961), .CP(clk), .RN(rst_n), .Q(y_z2[9])
         );
  HS65_GS_DFPRQX4 \data_out_reg[8]  ( .D(n1962), .CP(clk), .RN(rst_n), .Q(
        data_out[8]) );
  HS65_GS_DFPRQX4 \y_z1_reg[8]  ( .D(n1963), .CP(clk), .RN(rst_n), .Q(y_z1[8])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[8]  ( .D(n1964), .CP(clk), .RN(rst_n), .Q(y_z2[8])
         );
  HS65_GS_DFPRQX4 \data_out_reg[7]  ( .D(n1965), .CP(clk), .RN(rst_n), .Q(
        data_out[7]) );
  HS65_GS_DFPRQX4 \y_z1_reg[7]  ( .D(n1966), .CP(clk), .RN(rst_n), .Q(y_z1[7])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[7]  ( .D(n1967), .CP(clk), .RN(rst_n), .Q(y_z2[7])
         );
  HS65_GS_DFPRQX4 \data_out_reg[6]  ( .D(n1968), .CP(clk), .RN(rst_n), .Q(
        data_out[6]) );
  HS65_GS_DFPRQX4 \y_z1_reg[6]  ( .D(n1969), .CP(clk), .RN(rst_n), .Q(y_z1[6])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[6]  ( .D(n1970), .CP(clk), .RN(rst_n), .Q(y_z2[6])
         );
  HS65_GS_DFPRQX4 \data_out_reg[5]  ( .D(n1971), .CP(clk), .RN(rst_n), .Q(
        data_out[5]) );
  HS65_GS_DFPRQX4 \y_z1_reg[5]  ( .D(n1972), .CP(clk), .RN(rst_n), .Q(y_z1[5])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[5]  ( .D(n1973), .CP(clk), .RN(rst_n), .Q(y_z2[5])
         );
  HS65_GS_DFPRQX4 \data_out_reg[4]  ( .D(n1974), .CP(clk), .RN(rst_n), .Q(
        data_out[4]) );
  HS65_GS_DFPRQX4 \y_z1_reg[4]  ( .D(n1975), .CP(clk), .RN(rst_n), .Q(y_z1[4])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[4]  ( .D(n1976), .CP(clk), .RN(rst_n), .Q(y_z2[4])
         );
  HS65_GS_DFPRQX4 \data_out_reg[3]  ( .D(n1977), .CP(clk), .RN(rst_n), .Q(
        data_out[3]) );
  HS65_GS_DFPRQX4 \y_z1_reg[3]  ( .D(n1978), .CP(clk), .RN(rst_n), .Q(y_z1[3])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[3]  ( .D(n1979), .CP(clk), .RN(rst_n), .Q(y_z2[3])
         );
  HS65_GS_DFPRQX4 \data_out_reg[2]  ( .D(n1980), .CP(clk), .RN(rst_n), .Q(
        data_out[2]) );
  HS65_GS_DFPRQX4 \y_z1_reg[2]  ( .D(n1981), .CP(clk), .RN(rst_n), .Q(y_z1[2])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[2]  ( .D(n1982), .CP(clk), .RN(rst_n), .Q(y_z2[2])
         );
  HS65_GS_DFPRQX4 \data_out_reg[1]  ( .D(n1983), .CP(clk), .RN(rst_n), .Q(
        data_out[1]) );
  HS65_GS_DFPRQX4 \y_z1_reg[1]  ( .D(n1984), .CP(clk), .RN(rst_n), .Q(y_z1[1])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[1]  ( .D(n1985), .CP(clk), .RN(rst_n), .Q(
        \mul_a2/fa1_s0[1] ) );
  HS65_GS_DFPRQX4 \data_out_reg[0]  ( .D(n1986), .CP(clk), .RN(rst_n), .Q(
        data_out[0]) );
  HS65_GS_DFPRQX4 \y_z1_reg[0]  ( .D(n1987), .CP(clk), .RN(rst_n), .Q(y_z1[0])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[0]  ( .D(n1988), .CP(clk), .RN(rst_n), .Q(
        \mul_a2/fa1_s0[0] ) );
  HS65_GS_NOR2X3 U3 ( .A(y_z2[15]), .B(n1287), .Z(n1) );
  HS65_GS_NOR2X3 U4 ( .A(y_z2[15]), .B(n1224), .Z(n2) );
  HS65_GS_AND2X4 U5 ( .A(\mul_b1/fa1_s1_r[32] ), .B(\mul_b1/fa1_s0_r[32] ), 
        .Z(n222) );
  HS65_GSS_XOR2X3 U6 ( .A(\mul_b1/fa1_s0_r[31] ), .B(\mul_b1/fa1_s1_r[31] ), 
        .Z(n213) );
  HS65_GS_AND2X4 U7 ( .A(\mul_b1/fa1_s1_r[30] ), .B(\mul_b1/fa1_s0_r[30] ), 
        .Z(n212) );
  HS65_GSS_XOR2X3 U8 ( .A(\mul_b1/fa1_s0_r[32] ), .B(\mul_b1/fa1_s1_r[32] ), 
        .Z(n4) );
  HS65_GS_AND2X4 U9 ( .A(\mul_b1/fa1_s1_r[31] ), .B(\mul_b1/fa1_s0_r[31] ), 
        .Z(n3) );
  HS65_GS_AND2X4 U10 ( .A(n215), .B(n214), .Z(n6) );
  HS65_GS_FA1X4 U11 ( .A0(n4), .B0(\mul_b1/fa1_s2_r[32] ), .CI(n3), .CO(n5), 
        .S0(n214) );
  HS65_GSS_XOR2X3 U12 ( .A(n6), .B(n5), .Z(n219) );
  HS65_GS_AND2X4 U13 ( .A(\mul_b1/fa1_s0_r[27] ), .B(\mul_b1/fa1_s1_r[27] ), 
        .Z(n7) );
  HS65_GSS_XOR2X3 U14 ( .A(\mul_b1/fa1_s0_r[28] ), .B(\mul_b1/fa1_s1_r[28] ), 
        .Z(n18) );
  HS65_GS_NAND2X2 U15 ( .A(n19), .B(n18), .Z(n17) );
  HS65_GS_IVX2 U16 ( .A(n17), .Z(n11) );
  HS65_GS_FA1X4 U17 ( .A0(\mul_b1/fa1_c2_r[27] ), .B0(\mul_b1/fa1_s2_r[28] ), 
        .CI(n7), .CO(n12), .S0(n19) );
  HS65_GS_NOR2X2 U18 ( .A(n11), .B(n12), .Z(n13) );
  HS65_GS_AND2X4 U19 ( .A(\mul_b1/fa1_s1_r[28] ), .B(\mul_b1/fa1_s0_r[28] ), 
        .Z(n205) );
  HS65_GS_NAND2X2 U20 ( .A(\mul_b1/fa1_s2_r[29] ), .B(\mul_b1/fa1_c2_r[28] ), 
        .Z(n199) );
  HS65_GS_OA12X4 U21 ( .A(\mul_b1/fa1_s2_r[29] ), .B(\mul_b1/fa1_c2_r[28] ), 
        .C(n199), .Z(n8) );
  HS65_GS_AND2X4 U22 ( .A(n205), .B(n8), .Z(n202) );
  HS65_GSS_XOR2X3 U23 ( .A(\mul_b1/fa1_s0_r[29] ), .B(\mul_b1/fa1_s1_r[29] ), 
        .Z(n203) );
  HS65_GS_NOR2X2 U24 ( .A(n205), .B(n8), .Z(n200) );
  HS65_GS_OAI21X2 U25 ( .A(n202), .B(n200), .C(n203), .Z(n9) );
  HS65_GS_OAI13X1 U26 ( .A(n202), .B(n203), .C(n200), .D(n9), .Z(n198) );
  HS65_GS_NAND3X2 U27 ( .A(\mul_b1/fa1_c2_r[27] ), .B(\mul_b1/fa1_s2_r[28] ), 
        .C(n11), .Z(n10) );
  HS65_GS_OAI21X2 U28 ( .A(n12), .B(n11), .C(n10), .Z(n197) );
  HS65_GS_NOR2X2 U29 ( .A(n198), .B(n197), .Z(n196) );
  HS65_GS_NOR2X2 U30 ( .A(n13), .B(n196), .Z(n1011) );
  HS65_GS_AND2X4 U31 ( .A(\mul_b1/fa1_s0_r[26] ), .B(\mul_b1/fa1_s1_r[26] ), 
        .Z(n14) );
  HS65_GSS_XOR2X3 U32 ( .A(\mul_b1/fa1_s0_r[27] ), .B(\mul_b1/fa1_s1_r[27] ), 
        .Z(n25) );
  HS65_GS_NAND2X2 U33 ( .A(n26), .B(n25), .Z(n24) );
  HS65_GS_IVX2 U34 ( .A(n24), .Z(n16) );
  HS65_GS_FA1X4 U35 ( .A0(\mul_b1/fa1_c2_r[26] ), .B0(\mul_b1/fa1_s2_r[27] ), 
        .CI(n14), .CO(n15), .S0(n26) );
  HS65_GS_AOI12X2 U36 ( .A(n25), .B(n26), .C(n15), .Z(n20) );
  HS65_GS_AOI13X2 U37 ( .A(n16), .B(\mul_b1/fa1_s2_r[27] ), .C(
        \mul_b1/fa1_c2_r[26] ), .D(n20), .Z(n194) );
  HS65_GS_OAI21X2 U38 ( .A(n19), .B(n18), .C(n17), .Z(n193) );
  HS65_GS_AOI12X2 U39 ( .A(n194), .B(n193), .C(n20), .Z(n1005) );
  HS65_GSS_XOR2X3 U40 ( .A(\mul_b1/fa1_s0_r[26] ), .B(\mul_b1/fa1_s1_r[26] ), 
        .Z(n41) );
  HS65_GS_AND2X4 U41 ( .A(\mul_b1/fa1_s0_r[25] ), .B(\mul_b1/fa1_s1_r[25] ), 
        .Z(n21) );
  HS65_GS_FA1X4 U42 ( .A0(\mul_b1/fa1_c2_r[25] ), .B0(\mul_b1/fa1_s2_r[26] ), 
        .CI(n21), .CO(n22), .S0(n42) );
  HS65_GS_AOI12X2 U43 ( .A(n41), .B(n42), .C(n22), .Z(n28) );
  HS65_GS_NAND2X2 U44 ( .A(n42), .B(n41), .Z(n40) );
  HS65_GS_IVX2 U45 ( .A(n40), .Z(n23) );
  HS65_GS_AOI13X2 U46 ( .A(n23), .B(\mul_b1/fa1_s2_r[26] ), .C(
        \mul_b1/fa1_c2_r[25] ), .D(n28), .Z(n30) );
  HS65_GS_OAI21X2 U47 ( .A(n26), .B(n25), .C(n24), .Z(n29) );
  HS65_GS_AND2X4 U48 ( .A(n30), .B(n29), .Z(n27) );
  HS65_GS_NOR2X2 U49 ( .A(n28), .B(n27), .Z(n192) );
  HS65_GSS_XOR2X3 U50 ( .A(n30), .B(n29), .Z(n1019) );
  HS65_GS_AND2X4 U51 ( .A(\mul_b1/fa1_s0_r[23] ), .B(\mul_b1/fa1_s1_r[23] ), 
        .Z(n31) );
  HS65_GSS_XOR2X3 U52 ( .A(\mul_b1/fa1_s0_r[24] ), .B(\mul_b1/fa1_s1_r[24] ), 
        .Z(n49) );
  HS65_GS_NAND2X2 U53 ( .A(n50), .B(n49), .Z(n48) );
  HS65_GS_IVX2 U54 ( .A(n48), .Z(n33) );
  HS65_GS_FA1X4 U55 ( .A0(\mul_b1/fa1_c2_r[23] ), .B0(\mul_b1/fa1_s2_r[24] ), 
        .CI(n31), .CO(n32), .S0(n50) );
  HS65_GS_AOI12X2 U56 ( .A(n49), .B(n50), .C(n32), .Z(n34) );
  HS65_GS_AOI13X2 U57 ( .A(n33), .B(\mul_b1/fa1_c2_r[23] ), .C(
        \mul_b1/fa1_s2_r[24] ), .D(n34), .Z(n187) );
  HS65_GS_AND2X4 U58 ( .A(\mul_b1/fa1_s0_r[24] ), .B(\mul_b1/fa1_s1_r[24] ), 
        .Z(n36) );
  HS65_GSS_XOR2X3 U59 ( .A(\mul_b1/fa1_s0_r[25] ), .B(\mul_b1/fa1_s1_r[25] ), 
        .Z(n38) );
  HS65_GS_NAND2X2 U60 ( .A(n37), .B(n38), .Z(n35) );
  HS65_GS_OAI21X2 U61 ( .A(n37), .B(n38), .C(n35), .Z(n186) );
  HS65_GS_NAND2X2 U62 ( .A(n187), .B(n186), .Z(n185) );
  HS65_GS_NOR2AX3 U63 ( .A(n185), .B(n34), .Z(n1442) );
  HS65_GS_IVX2 U64 ( .A(n35), .Z(n190) );
  HS65_GS_FA1X4 U65 ( .A0(\mul_b1/fa1_c2_r[24] ), .B0(\mul_b1/fa1_s2_r[25] ), 
        .CI(n36), .CO(n189), .S0(n37) );
  HS65_GS_AOI12X2 U66 ( .A(n38), .B(n37), .C(n189), .Z(n39) );
  HS65_GS_AOI13X2 U67 ( .A(n190), .B(\mul_b1/fa1_s2_r[25] ), .C(
        \mul_b1/fa1_c2_r[24] ), .D(n39), .Z(n44) );
  HS65_GS_OAI21X2 U68 ( .A(n42), .B(n41), .C(n40), .Z(n43) );
  HS65_GS_NAND2X2 U69 ( .A(n44), .B(n43), .Z(n188) );
  HS65_GS_OAI21X2 U70 ( .A(n44), .B(n43), .C(n188), .Z(n1441) );
  HS65_GS_AND2X4 U71 ( .A(\mul_b1/fa1_s0_r[22] ), .B(\mul_b1/fa1_s1_r[22] ), 
        .Z(n45) );
  HS65_GSS_XOR2X3 U72 ( .A(\mul_b1/fa1_s0_r[23] ), .B(\mul_b1/fa1_s1_r[23] ), 
        .Z(n56) );
  HS65_GS_NAND2X2 U73 ( .A(n57), .B(n56), .Z(n55) );
  HS65_GS_IVX2 U74 ( .A(n55), .Z(n47) );
  HS65_GS_FA1X4 U75 ( .A0(\mul_b1/fa1_c2_r[22] ), .B0(\mul_b1/fa1_s2_r[23] ), 
        .CI(n45), .CO(n46), .S0(n57) );
  HS65_GS_AOI12X2 U76 ( .A(n56), .B(n57), .C(n46), .Z(n51) );
  HS65_GS_AOI13X2 U77 ( .A(n47), .B(\mul_b1/fa1_c2_r[22] ), .C(
        \mul_b1/fa1_s2_r[23] ), .D(n51), .Z(n184) );
  HS65_GS_OAI21X2 U78 ( .A(n50), .B(n49), .C(n48), .Z(n183) );
  HS65_GS_NAND2X2 U79 ( .A(n184), .B(n183), .Z(n182) );
  HS65_GS_NOR2AX3 U80 ( .A(n182), .B(n51), .Z(n1446) );
  HS65_GS_AND2X4 U81 ( .A(\mul_b1/fa1_s0_r[21] ), .B(\mul_b1/fa1_s1_r[21] ), 
        .Z(n52) );
  HS65_GSS_XOR2X3 U82 ( .A(\mul_b1/fa1_s0_r[22] ), .B(\mul_b1/fa1_s1_r[22] ), 
        .Z(n173) );
  HS65_GS_NAND2X2 U83 ( .A(n174), .B(n173), .Z(n172) );
  HS65_GS_IVX2 U84 ( .A(n172), .Z(n54) );
  HS65_GS_FA1X4 U85 ( .A0(\mul_b1/fa1_c2_r[21] ), .B0(\mul_b1/fa1_s2_r[22] ), 
        .CI(n52), .CO(n53), .S0(n174) );
  HS65_GS_AOI12X2 U86 ( .A(n173), .B(n174), .C(n53), .Z(n58) );
  HS65_GS_AOI13X2 U87 ( .A(n54), .B(\mul_b1/fa1_c2_r[21] ), .C(
        \mul_b1/fa1_s2_r[22] ), .D(n58), .Z(n181) );
  HS65_GS_OAI21X2 U88 ( .A(n57), .B(n56), .C(n55), .Z(n180) );
  HS65_GS_NAND2X2 U89 ( .A(n181), .B(n180), .Z(n179) );
  HS65_GS_NOR2AX3 U90 ( .A(n179), .B(n58), .Z(n1450) );
  HS65_GS_NAND2X2 U91 ( .A(n68), .B(n67), .Z(n66) );
  HS65_GS_IVX2 U92 ( .A(n66), .Z(n61) );
  HS65_GS_FA1X4 U93 ( .A0(\mul_b1/fa1_c2_r[19] ), .B0(\mul_b1/fa1_s2_r[20] ), 
        .CI(n59), .CO(n60), .S0(n68) );
  HS65_GS_AOI12X2 U94 ( .A(n67), .B(n68), .C(n60), .Z(n62) );
  HS65_GS_AOI13X2 U95 ( .A(n61), .B(\mul_b1/fa1_c2_r[19] ), .C(
        \mul_b1/fa1_s2_r[20] ), .D(n62), .Z(n165) );
  HS65_GS_FA1X4 U96 ( .A0(\mul_b1/fa1_s0_r[20] ), .B0(\mul_b1/fa1_s1_r[20] ), 
        .CI(\mul_b1/fa1_c0_r[19] ), .CO(n167), .S0(n67) );
  HS65_GSS_XOR2X3 U97 ( .A(\mul_b1/fa1_s0_r[21] ), .B(\mul_b1/fa1_s1_r[21] ), 
        .Z(n170) );
  HS65_GS_NAND2X2 U98 ( .A(n169), .B(n170), .Z(n166) );
  HS65_GS_OAI21X2 U99 ( .A(n169), .B(n170), .C(n166), .Z(n164) );
  HS65_GS_NAND2X2 U100 ( .A(n165), .B(n164), .Z(n163) );
  HS65_GS_NOR2AX3 U101 ( .A(n163), .B(n62), .Z(n1458) );
  HS65_GS_FA1X4 U102 ( .A0(\mul_b1/fa1_s0_r[19] ), .B0(\mul_b1/fa1_s1_r[19] ), 
        .CI(\mul_b1/fa1_c0_r[18] ), .CO(n59), .S0(n154) );
  HS65_GS_NAND2X2 U103 ( .A(n155), .B(n154), .Z(n153) );
  HS65_GS_IVX2 U104 ( .A(n153), .Z(n65) );
  HS65_GS_FA1X4 U105 ( .A0(\mul_b1/fa1_c2_r[18] ), .B0(\mul_b1/fa1_s2_r[19] ), 
        .CI(n63), .CO(n64), .S0(n155) );
  HS65_GS_AOI12X2 U106 ( .A(n154), .B(n155), .C(n64), .Z(n69) );
  HS65_GS_AOI13X2 U107 ( .A(n65), .B(\mul_b1/fa1_c2_r[18] ), .C(
        \mul_b1/fa1_s2_r[19] ), .D(n69), .Z(n162) );
  HS65_GS_OAI21X2 U108 ( .A(n68), .B(n67), .C(n66), .Z(n161) );
  HS65_GS_NAND2X2 U109 ( .A(n162), .B(n161), .Z(n160) );
  HS65_GS_NOR2AX3 U110 ( .A(n160), .B(n69), .Z(n1462) );
  HS65_GS_NAND2X2 U111 ( .A(n79), .B(n78), .Z(n77) );
  HS65_GS_IVX2 U112 ( .A(n77), .Z(n72) );
  HS65_GS_FA1X4 U113 ( .A0(\mul_b1/fa1_c2_r[16] ), .B0(\mul_b1/fa1_s2_r[17] ), 
        .CI(n70), .CO(n71), .S0(n79) );
  HS65_GS_AOI12X2 U114 ( .A(n78), .B(n79), .C(n71), .Z(n73) );
  HS65_GS_AOI13X2 U115 ( .A(n72), .B(\mul_b1/fa1_c2_r[16] ), .C(
        \mul_b1/fa1_s2_r[17] ), .D(n73), .Z(n146) );
  HS65_GS_FA1X4 U116 ( .A0(\mul_b1/fa1_s0_r[17] ), .B0(\mul_b1/fa1_s1_r[17] ), 
        .CI(\mul_b1/fa1_c0_r[16] ), .CO(n148), .S0(n78) );
  HS65_GS_FA1X4 U117 ( .A0(\mul_b1/fa1_s0_r[18] ), .B0(\mul_b1/fa1_s1_r[18] ), 
        .CI(\mul_b1/fa1_c0_r[17] ), .CO(n63), .S0(n151) );
  HS65_GS_NAND2X2 U118 ( .A(n150), .B(n151), .Z(n147) );
  HS65_GS_OAI21X2 U119 ( .A(n150), .B(n151), .C(n147), .Z(n145) );
  HS65_GS_NAND2X2 U120 ( .A(n146), .B(n145), .Z(n144) );
  HS65_GS_NOR2AX3 U121 ( .A(n144), .B(n73), .Z(n1470) );
  HS65_GS_FA1X4 U122 ( .A0(\mul_b1/fa1_s0_r[16] ), .B0(\mul_b1/fa1_s1_r[16] ), 
        .CI(\mul_b1/fa1_c0_r[15] ), .CO(n70), .S0(n85) );
  HS65_GS_NAND2X2 U123 ( .A(n86), .B(n85), .Z(n84) );
  HS65_GS_IVX2 U124 ( .A(n84), .Z(n76) );
  HS65_GS_FA1X4 U125 ( .A0(\mul_b1/fa1_c2_r[15] ), .B0(\mul_b1/fa1_s2_r[16] ), 
        .CI(n74), .CO(n75), .S0(n86) );
  HS65_GS_NOR2X2 U126 ( .A(n76), .B(n75), .Z(n80) );
  HS65_GS_AOI13X2 U127 ( .A(n76), .B(\mul_b1/fa1_c2_r[15] ), .C(
        \mul_b1/fa1_s2_r[16] ), .D(n80), .Z(n143) );
  HS65_GS_OAI21X2 U128 ( .A(n79), .B(n78), .C(n77), .Z(n142) );
  HS65_GS_NAND2X2 U129 ( .A(n143), .B(n142), .Z(n141) );
  HS65_GS_NOR2AX3 U130 ( .A(n141), .B(n80), .Z(n1474) );
  HS65_GS_FA1X4 U131 ( .A0(\mul_b1/fa1_s0_r[15] ), .B0(\mul_b1/fa1_s1_r[15] ), 
        .CI(\mul_b1/fa1_c0_r[14] ), .CO(n74), .S0(n81) );
  HS65_GS_AND2X4 U132 ( .A(n92), .B(n91), .Z(n83) );
  HS65_GS_FA1X4 U133 ( .A0(\mul_b1/fa1_c2_r[14] ), .B0(\mul_b1/fa1_s2_r[15] ), 
        .CI(n81), .CO(n82), .S0(n92) );
  HS65_GS_AOI12X2 U134 ( .A(n91), .B(n92), .C(n82), .Z(n87) );
  HS65_GS_AOI13X2 U135 ( .A(n83), .B(\mul_b1/fa1_s2_r[15] ), .C(
        \mul_b1/fa1_c2_r[14] ), .D(n87), .Z(n89) );
  HS65_GS_OAI21X2 U136 ( .A(n86), .B(n85), .C(n84), .Z(n88) );
  HS65_GS_AOI12X2 U137 ( .A(n89), .B(n88), .C(n87), .Z(n1477) );
  HS65_GSS_XOR2X3 U138 ( .A(n89), .B(n88), .Z(n1480) );
  HS65_GS_PAO2X4 U139 ( .A(\mul_b1/fa1_c0_r[12] ), .B(\mul_b1/fa1_s1_r[13] ), 
        .P(\mul_b1/fa1_s0_r[13] ), .Z(n94) );
  HS65_GS_FA1X4 U140 ( .A0(\mul_b1/fa1_s0_r[14] ), .B0(\mul_b1/fa1_s1_r[14] ), 
        .CI(\mul_b1/fa1_c0_r[13] ), .CO(n91), .S0(n93) );
  HS65_GS_PAOI2X1 U141 ( .A(\mul_b1/fa1_c0_r[11] ), .B(\mul_b1/fa1_s1_r[12] ), 
        .P(\mul_b1/fa1_s0_r[12] ), .Z(n96) );
  HS65_GSS_XNOR3X2 U142 ( .A(\mul_b1/fa1_c0_r[12] ), .B(\mul_b1/fa1_s1_r[13] ), 
        .C(\mul_b1/fa1_s0_r[13] ), .Z(n95) );
  HS65_GS_IVX2 U143 ( .A(\mul_b1/fa1_s2_r[13] ), .Z(n90) );
  HS65_GS_PAOI2X1 U144 ( .A(n96), .B(n95), .P(n90), .Z(n135) );
  HS65_GS_NAND2X2 U145 ( .A(n136), .B(n135), .Z(n134) );
  HS65_GS_IVX2 U146 ( .A(n134), .Z(n139) );
  HS65_GSS_XOR2X3 U147 ( .A(n92), .B(n91), .Z(n138) );
  HS65_GS_FA1X4 U148 ( .A0(\mul_b1/fa1_s2_r[14] ), .B0(n94), .CI(n93), .CO(
        n137), .S0(n136) );
  HS65_GSS_XNOR3X2 U149 ( .A(\mul_b1/fa1_c0_r[11] ), .B(\mul_b1/fa1_s1_r[12] ), 
        .C(\mul_b1/fa1_s0_r[12] ), .Z(n97) );
  HS65_GS_PAOI2X1 U150 ( .A(\mul_b1/fa1_c0_r[10] ), .B(\mul_b1/fa1_s1_r[11] ), 
        .P(\mul_b1/fa1_s0_r[11] ), .Z(n98) );
  HS65_GS_NOR2X2 U151 ( .A(n97), .B(n98), .Z(n133) );
  HS65_GSS_XOR3X2 U152 ( .A(n96), .B(\mul_b1/fa1_s2_r[13] ), .C(n95), .Z(n132)
         );
  HS65_GS_IVX2 U153 ( .A(n132), .Z(n130) );
  HS65_GSS_XNOR3X2 U154 ( .A(\mul_b1/fa1_c0_r[10] ), .B(\mul_b1/fa1_s1_r[11] ), 
        .C(\mul_b1/fa1_s0_r[11] ), .Z(n119) );
  HS65_GS_PAOI2X1 U155 ( .A(\mul_b1/fa1_s1_r[10] ), .B(\mul_b1/fa1_c0_r[9] ), 
        .P(\mul_b1/fa1_s0_r[10] ), .Z(n120) );
  HS65_GS_NOR2X2 U156 ( .A(n119), .B(n120), .Z(n128) );
  HS65_GSS_XOR2X3 U157 ( .A(n98), .B(n97), .Z(n127) );
  HS65_GSS_XNOR3X2 U158 ( .A(\mul_b1/fa1_c0_r[8] ), .B(\mul_b1/fa1_s1_r[9] ), 
        .C(\mul_b1/fa1_s0_r[9] ), .Z(n110) );
  HS65_GS_NAND2X2 U159 ( .A(\mul_b1/fa1_c0_r[7] ), .B(\mul_b1/fa1_s0_r[8] ), 
        .Z(n99) );
  HS65_GS_NOR2X2 U160 ( .A(n110), .B(n99), .Z(n118) );
  HS65_GS_PAOI2X1 U161 ( .A(\mul_b1/fa1_c0_r[8] ), .B(\mul_b1/fa1_s1_r[9] ), 
        .P(\mul_b1/fa1_s0_r[9] ), .Z(n121) );
  HS65_GSS_XNOR3X2 U162 ( .A(\mul_b1/fa1_s1_r[10] ), .B(\mul_b1/fa1_c0_r[9] ), 
        .C(\mul_b1/fa1_s0_r[10] ), .Z(n122) );
  HS65_GSS_XOR2X3 U163 ( .A(n121), .B(n122), .Z(n117) );
  HS65_GS_NAND2X2 U164 ( .A(\mul_b1/fa1_c0_r[5] ), .B(\mul_b1/fa1_s0_r[6] ), 
        .Z(n100) );
  HS65_GSS_XNOR2X3 U165 ( .A(\mul_b1/fa1_c0_r[6] ), .B(\mul_b1/fa1_s0_r[7] ), 
        .Z(n101) );
  HS65_GS_NOR2X2 U166 ( .A(n100), .B(n101), .Z(n109) );
  HS65_GSS_XNOR2X3 U167 ( .A(\mul_b1/fa1_c0_r[7] ), .B(\mul_b1/fa1_s0_r[8] ), 
        .Z(n111) );
  HS65_GS_IVX2 U168 ( .A(n111), .Z(n108) );
  HS65_GS_IVX2 U169 ( .A(n101), .Z(n105) );
  HS65_GS_NAND2X2 U170 ( .A(\mul_b1/fa1_c0_r[4] ), .B(\mul_b1/fa1_s0_r[5] ), 
        .Z(n103) );
  HS65_GSS_XNOR2X3 U171 ( .A(\mul_b1/fa1_c0_r[5] ), .B(\mul_b1/fa1_s0_r[6] ), 
        .Z(n102) );
  HS65_GS_NOR2X2 U172 ( .A(n103), .B(n102), .Z(n104) );
  HS65_GS_NAND2X2 U173 ( .A(n105), .B(n104), .Z(n106) );
  HS65_GS_NOR2X2 U174 ( .A(n111), .B(n106), .Z(n107) );
  HS65_GS_AO12X4 U175 ( .A(n109), .B(n108), .C(n107), .Z(n115) );
  HS65_GS_IVX2 U176 ( .A(n110), .Z(n114) );
  HS65_GS_NAND2X2 U177 ( .A(\mul_b1/fa1_c0_r[6] ), .B(\mul_b1/fa1_s0_r[7] ), 
        .Z(n112) );
  HS65_GS_NOR2X2 U178 ( .A(n112), .B(n111), .Z(n113) );
  HS65_GS_PAO2X4 U179 ( .A(n115), .B(n114), .P(n113), .Z(n116) );
  HS65_GS_PAO2X4 U180 ( .A(n118), .B(n117), .P(n116), .Z(n125) );
  HS65_GSS_XOR2X3 U181 ( .A(n120), .B(n119), .Z(n124) );
  HS65_GS_NOR2X2 U182 ( .A(n122), .B(n121), .Z(n123) );
  HS65_GS_PAO2X4 U183 ( .A(n125), .B(n124), .P(n123), .Z(n126) );
  HS65_GS_PAOI2X1 U184 ( .A(n128), .B(n127), .P(n126), .Z(n129) );
  HS65_GS_NOR2X2 U185 ( .A(n130), .B(n129), .Z(n131) );
  HS65_GS_AOI12X2 U186 ( .A(n133), .B(n132), .C(n131), .Z(n1872) );
  HS65_GS_OAI21X2 U187 ( .A(n136), .B(n135), .C(n134), .Z(n1871) );
  HS65_GS_NOR2X2 U188 ( .A(n1872), .B(n1871), .Z(n1870) );
  HS65_GS_AND2X4 U189 ( .A(n1484), .B(n1870), .Z(n1486) );
  HS65_GS_FA1X4 U190 ( .A0(n139), .B0(n138), .CI(n137), .CO(n140), .S0(n1484)
         );
  HS65_GS_NOR2X2 U191 ( .A(n1486), .B(n140), .Z(n1481) );
  HS65_GS_NOR2X2 U192 ( .A(n1480), .B(n1481), .Z(n1479) );
  HS65_GS_OAI21X2 U193 ( .A(n143), .B(n142), .C(n141), .Z(n1476) );
  HS65_GS_OAI21X2 U194 ( .A(n146), .B(n145), .C(n144), .Z(n1472) );
  HS65_GS_IVX2 U195 ( .A(n147), .Z(n152) );
  HS65_GS_FA1X4 U196 ( .A0(\mul_b1/fa1_c2_r[17] ), .B0(\mul_b1/fa1_s2_r[18] ), 
        .CI(n148), .CO(n149), .S0(n150) );
  HS65_GS_AOI12X2 U197 ( .A(n151), .B(n150), .C(n149), .Z(n158) );
  HS65_GS_AOI13X2 U198 ( .A(n152), .B(\mul_b1/fa1_c2_r[17] ), .C(
        \mul_b1/fa1_s2_r[18] ), .D(n158), .Z(n157) );
  HS65_GS_OAI21X2 U199 ( .A(n155), .B(n154), .C(n153), .Z(n156) );
  HS65_GS_NAND2X2 U200 ( .A(n157), .B(n156), .Z(n159) );
  HS65_GS_OAI21X2 U201 ( .A(n157), .B(n156), .C(n159), .Z(n1468) );
  HS65_GS_NOR2AX3 U202 ( .A(n159), .B(n158), .Z(n1465) );
  HS65_GS_OAI21X2 U203 ( .A(n162), .B(n161), .C(n160), .Z(n1464) );
  HS65_GS_OAI21X2 U204 ( .A(n165), .B(n164), .C(n163), .Z(n1460) );
  HS65_GS_IVX2 U205 ( .A(n166), .Z(n171) );
  HS65_GS_FA1X4 U206 ( .A0(\mul_b1/fa1_c2_r[20] ), .B0(\mul_b1/fa1_s2_r[21] ), 
        .CI(n167), .CO(n168), .S0(n169) );
  HS65_GS_AOI12X2 U207 ( .A(n170), .B(n169), .C(n168), .Z(n177) );
  HS65_GS_AOI13X2 U208 ( .A(n171), .B(\mul_b1/fa1_c2_r[20] ), .C(
        \mul_b1/fa1_s2_r[21] ), .D(n177), .Z(n176) );
  HS65_GS_OAI21X2 U209 ( .A(n174), .B(n173), .C(n172), .Z(n175) );
  HS65_GS_NAND2X2 U210 ( .A(n176), .B(n175), .Z(n178) );
  HS65_GS_OAI21X2 U211 ( .A(n176), .B(n175), .C(n178), .Z(n1456) );
  HS65_GS_NOR2AX3 U212 ( .A(n178), .B(n177), .Z(n1453) );
  HS65_GS_OAI21X2 U213 ( .A(n181), .B(n180), .C(n179), .Z(n1452) );
  HS65_GS_OAI21X2 U214 ( .A(n184), .B(n183), .C(n182), .Z(n1448) );
  HS65_GS_OAI21X2 U215 ( .A(n187), .B(n186), .C(n185), .Z(n1444) );
  HS65_GS_IVX2 U216 ( .A(n997), .Z(n998) );
  HS65_GS_OAI21X2 U217 ( .A(n190), .B(n189), .C(n188), .Z(n996) );
  HS65_GS_PAOI2X1 U218 ( .A(n1019), .B(n998), .P(n996), .Z(n191) );
  HS65_GS_NOR2X2 U219 ( .A(n192), .B(n191), .Z(n1875) );
  HS65_GS_AND2X4 U220 ( .A(n192), .B(n191), .Z(n1874) );
  HS65_GSS_XNOR2X3 U221 ( .A(n194), .B(n193), .Z(n1877) );
  HS65_GS_NOR2X2 U222 ( .A(n1874), .B(n1877), .Z(n195) );
  HS65_GS_NOR2X2 U223 ( .A(n1875), .B(n195), .Z(n1004) );
  HS65_GS_AO12X4 U224 ( .A(n198), .B(n197), .C(n196), .Z(n1003) );
  HS65_GS_AND2X4 U225 ( .A(\mul_b1/fa1_s1_r[29] ), .B(\mul_b1/fa1_s0_r[29] ), 
        .Z(n211) );
  HS65_GSS_XOR2X3 U226 ( .A(\mul_b1/fa1_s0_r[30] ), .B(\mul_b1/fa1_s1_r[30] ), 
        .Z(n210) );
  HS65_GS_IVX2 U227 ( .A(n199), .Z(n204) );
  HS65_GS_NOR2AX3 U228 ( .A(n203), .B(n200), .Z(n201) );
  HS65_GS_NOR3X1 U229 ( .A(n204), .B(n202), .C(n201), .Z(n209) );
  HS65_GS_AO31X4 U230 ( .A(n205), .B(n204), .C(n203), .D(n209), .Z(n206) );
  HS65_GS_NOR2X2 U231 ( .A(n207), .B(n206), .Z(n208) );
  HS65_GS_AO12X4 U232 ( .A(n207), .B(n206), .C(n208), .Z(n1009) );
  HS65_GS_NOR2X2 U233 ( .A(n209), .B(n208), .Z(n1000) );
  HS65_GS_FA1X4 U234 ( .A0(n211), .B0(n210), .CI(\mul_b1/fa1_s2_r[30] ), .CO(
        n217), .S0(n207) );
  HS65_GS_FA1X4 U235 ( .A0(\mul_b1/fa1_s2_r[31] ), .B0(n213), .CI(n212), .CO(
        n215), .S0(n216) );
  HS65_GSS_XOR2X3 U236 ( .A(n217), .B(n216), .Z(n999) );
  HS65_GSS_XOR2X3 U237 ( .A(n215), .B(n214), .Z(n1007) );
  HS65_GS_AND2X4 U238 ( .A(n217), .B(n216), .Z(n1006) );
  HS65_GSS_XOR2X3 U239 ( .A(n219), .B(n218), .Z(n220) );
  HS65_GSS_XOR3X2 U240 ( .A(\mul_b1/fa1_s0_r[33] ), .B(\mul_b1/fa1_s1_r[33] ), 
        .C(n220), .Z(n221) );
  HS65_GSS_XOR3X2 U241 ( .A(n222), .B(\mul_b1/fa1_s2_r[33] ), .C(n221), .Z(
        \mul_b1/result_sat[15] ) );
  HS65_GS_AND2X4 U242 ( .A(\mul_a2/fa1_c1_r[31] ), .B(\mul_a2/fa1_s2_r[32] ), 
        .Z(n423) );
  HS65_GSS_XOR2X3 U243 ( .A(\mul_a2/fa1_s2_r[31] ), .B(\mul_a2/fa1_c1_r[30] ), 
        .Z(n406) );
  HS65_GSS_XOR2X3 U244 ( .A(\mul_a2/fa1_s2_r[32] ), .B(\mul_a2/fa1_c1_r[31] ), 
        .Z(n415) );
  HS65_GS_FA1X4 U245 ( .A0(\mul_a2/fa1_s0_r[32] ), .B0(\mul_a2/fa1_s1_r[32] ), 
        .CI(\mul_a2/fa1_c0_r[31] ), .CO(n424), .S0(n414) );
  HS65_GS_FA1X4 U246 ( .A0(\mul_a2/fa1_s0_r[31] ), .B0(\mul_a2/fa1_s1_r[31] ), 
        .CI(\mul_a2/fa1_c0_r[30] ), .CO(n413), .S0(n405) );
  HS65_GS_AND2X4 U247 ( .A(\mul_a2/fa1_c1_r[30] ), .B(\mul_a2/fa1_s2_r[31] ), 
        .Z(n410) );
  HS65_GS_FA1X4 U248 ( .A0(\mul_a2/fa1_c1_r[28] ), .B0(\mul_a2/fa1_c2_r[28] ), 
        .CI(\mul_a2/fa1_s2_r[29] ), .CO(n400), .S0(n225) );
  HS65_GS_FA1X4 U249 ( .A0(\mul_a2/fa1_s0_r[29] ), .B0(\mul_a2/fa1_s1_r[29] ), 
        .CI(\mul_a2/fa1_c0_r[28] ), .CO(n403), .S0(n223) );
  HS65_GS_FA1X4 U250 ( .A0(\mul_a2/fa1_s0_r[30] ), .B0(\mul_a2/fa1_s1_r[30] ), 
        .CI(\mul_a2/fa1_c0_r[29] ), .CO(n404), .S0(n402) );
  HS65_GSS_XOR2X3 U251 ( .A(\mul_a2/fa1_s2_r[30] ), .B(\mul_a2/fa1_c1_r[29] ), 
        .Z(n401) );
  HS65_GS_FA1X4 U252 ( .A0(\mul_a2/fa1_c1_r[27] ), .B0(\mul_a2/fa1_c2_r[27] ), 
        .CI(\mul_a2/fa1_s2_r[28] ), .CO(n397), .S0(n228) );
  HS65_GS_FA1X4 U253 ( .A0(\mul_a2/fa1_s0_r[28] ), .B0(\mul_a2/fa1_s1_r[28] ), 
        .CI(\mul_a2/fa1_c0_r[27] ), .CO(n224), .S0(n226) );
  HS65_GS_FA1X4 U254 ( .A0(n225), .B0(n224), .CI(n223), .CO(n399), .S0(n395)
         );
  HS65_GS_FA1X4 U255 ( .A0(\mul_a2/fa1_c1_r[26] ), .B0(\mul_a2/fa1_c2_r[26] ), 
        .CI(\mul_a2/fa1_s2_r[27] ), .CO(n394), .S0(n388) );
  HS65_GS_FA1X4 U256 ( .A0(\mul_a2/fa1_s0_r[27] ), .B0(\mul_a2/fa1_s1_r[27] ), 
        .CI(\mul_a2/fa1_c0_r[26] ), .CO(n227), .S0(n386) );
  HS65_GS_FA1X4 U257 ( .A0(n228), .B0(n227), .CI(n226), .CO(n396), .S0(n392)
         );
  HS65_GS_FA1X4 U258 ( .A0(\mul_a2/fa1_c1_r[24] ), .B0(\mul_a2/fa1_c2_r[24] ), 
        .CI(\mul_a2/fa1_s2_r[25] ), .CO(n382), .S0(n231) );
  HS65_GS_FA1X4 U259 ( .A0(\mul_a2/fa1_s0_r[25] ), .B0(\mul_a2/fa1_s1_r[25] ), 
        .CI(\mul_a2/fa1_c0_r[24] ), .CO(n384), .S0(n229) );
  HS65_GS_FA1X4 U260 ( .A0(\mul_a2/fa1_s0_r[26] ), .B0(\mul_a2/fa1_s1_r[26] ), 
        .CI(\mul_a2/fa1_c0_r[25] ), .CO(n387), .S0(n383) );
  HS65_GS_FA1X4 U261 ( .A0(\mul_a2/fa1_c1_r[23] ), .B0(\mul_a2/fa1_c2_r[23] ), 
        .CI(\mul_a2/fa1_s2_r[24] ), .CO(n379), .S0(n234) );
  HS65_GS_FA1X4 U262 ( .A0(\mul_a2/fa1_s0_r[24] ), .B0(\mul_a2/fa1_s1_r[24] ), 
        .CI(\mul_a2/fa1_c0_r[23] ), .CO(n230), .S0(n232) );
  HS65_GS_FA1X4 U263 ( .A0(n231), .B0(n230), .CI(n229), .CO(n381), .S0(n377)
         );
  HS65_GS_FA1X4 U264 ( .A0(\mul_a2/fa1_c1_r[22] ), .B0(\mul_a2/fa1_c2_r[22] ), 
        .CI(\mul_a2/fa1_s2_r[23] ), .CO(n376), .S0(n370) );
  HS65_GS_FA1X4 U265 ( .A0(\mul_a2/fa1_s0_r[23] ), .B0(\mul_a2/fa1_s1_r[23] ), 
        .CI(\mul_a2/fa1_c0_r[22] ), .CO(n233), .S0(n368) );
  HS65_GS_FA1X4 U266 ( .A0(n234), .B0(n233), .CI(n232), .CO(n378), .S0(n374)
         );
  HS65_GS_FA1X4 U267 ( .A0(\mul_a2/fa1_c1_r[20] ), .B0(\mul_a2/fa1_c2_r[20] ), 
        .CI(\mul_a2/fa1_s2_r[21] ), .CO(n364), .S0(n237) );
  HS65_GS_FA1X4 U268 ( .A0(\mul_a2/fa1_s0_r[21] ), .B0(\mul_a2/fa1_s1_r[21] ), 
        .CI(\mul_a2/fa1_c0_r[20] ), .CO(n366), .S0(n235) );
  HS65_GS_FA1X4 U269 ( .A0(\mul_a2/fa1_s0_r[22] ), .B0(\mul_a2/fa1_s1_r[22] ), 
        .CI(\mul_a2/fa1_c0_r[21] ), .CO(n369), .S0(n365) );
  HS65_GS_FA1X4 U270 ( .A0(\mul_a2/fa1_c1_r[19] ), .B0(\mul_a2/fa1_c2_r[19] ), 
        .CI(\mul_a2/fa1_s2_r[20] ), .CO(n361), .S0(n240) );
  HS65_GS_FA1X4 U271 ( .A0(\mul_a2/fa1_s0_r[20] ), .B0(\mul_a2/fa1_s1_r[20] ), 
        .CI(\mul_a2/fa1_c0_r[19] ), .CO(n236), .S0(n238) );
  HS65_GS_FA1X4 U272 ( .A0(n237), .B0(n236), .CI(n235), .CO(n363), .S0(n359)
         );
  HS65_GS_FA1X4 U273 ( .A0(\mul_a2/fa1_c1_r[18] ), .B0(\mul_a2/fa1_c2_r[18] ), 
        .CI(\mul_a2/fa1_s2_r[19] ), .CO(n358), .S0(n243) );
  HS65_GS_FA1X4 U274 ( .A0(\mul_a2/fa1_s0_r[19] ), .B0(\mul_a2/fa1_s1_r[19] ), 
        .CI(\mul_a2/fa1_c0_r[18] ), .CO(n239), .S0(n241) );
  HS65_GS_FA1X4 U275 ( .A0(n240), .B0(n239), .CI(n238), .CO(n360), .S0(n356)
         );
  HS65_GS_FA1X4 U276 ( .A0(\mul_a2/fa1_c1_r[17] ), .B0(\mul_a2/fa1_c2_r[17] ), 
        .CI(\mul_a2/fa1_s2_r[18] ), .CO(n355), .S0(n246) );
  HS65_GS_FA1X4 U277 ( .A0(\mul_a2/fa1_s0_r[18] ), .B0(\mul_a2/fa1_s1_r[18] ), 
        .CI(\mul_a2/fa1_c0_r[17] ), .CO(n242), .S0(n244) );
  HS65_GS_FA1X4 U278 ( .A0(n243), .B0(n242), .CI(n241), .CO(n357), .S0(n353)
         );
  HS65_GS_FA1X4 U279 ( .A0(\mul_a2/fa1_c1_r[16] ), .B0(\mul_a2/fa1_c2_r[16] ), 
        .CI(\mul_a2/fa1_s2_r[17] ), .CO(n352), .S0(n249) );
  HS65_GS_FA1X4 U280 ( .A0(\mul_a2/fa1_s0_r[17] ), .B0(\mul_a2/fa1_s1_r[17] ), 
        .CI(\mul_a2/fa1_c0_r[16] ), .CO(n245), .S0(n247) );
  HS65_GS_FA1X4 U281 ( .A0(n246), .B0(n245), .CI(n244), .CO(n354), .S0(n350)
         );
  HS65_GS_FA1X4 U282 ( .A0(\mul_a2/fa1_c1_r[15] ), .B0(\mul_a2/fa1_c2_r[15] ), 
        .CI(\mul_a2/fa1_s2_r[16] ), .CO(n349), .S0(n252) );
  HS65_GS_FA1X4 U283 ( .A0(\mul_a2/fa1_s0_r[16] ), .B0(\mul_a2/fa1_s1_r[16] ), 
        .CI(\mul_a2/fa1_c0_r[15] ), .CO(n248), .S0(n250) );
  HS65_GS_FA1X4 U284 ( .A0(n249), .B0(n248), .CI(n247), .CO(n351), .S0(n347)
         );
  HS65_GS_FA1X4 U285 ( .A0(\mul_a2/fa1_s0_r[15] ), .B0(\mul_a2/fa1_s1_r[15] ), 
        .CI(\mul_a2/fa1_c0_r[14] ), .CO(n251), .S0(n255) );
  HS65_GS_FA1X4 U286 ( .A0(\mul_a2/fa1_c1_r[14] ), .B0(\mul_a2/fa1_c2_r[14] ), 
        .CI(\mul_a2/fa1_s2_r[15] ), .CO(n346), .S0(n254) );
  HS65_GS_FA1X4 U287 ( .A0(n252), .B0(n251), .CI(n250), .CO(n348), .S0(n344)
         );
  HS65_GS_AND2X4 U288 ( .A(\mul_a2/fa1_c1_r[13] ), .B(\mul_a2/fa1_s2_r[14] ), 
        .Z(n258) );
  HS65_GS_FA1X4 U289 ( .A0(n255), .B0(n254), .CI(n253), .CO(n345), .S0(n257)
         );
  HS65_GSS_XOR2X3 U290 ( .A(\mul_a2/fa1_c1_r[13] ), .B(\mul_a2/fa1_s2_r[14] ), 
        .Z(n337) );
  HS65_GS_FA1X4 U291 ( .A0(\mul_a2/fa1_s0_r[14] ), .B0(\mul_a2/fa1_s1_r[14] ), 
        .CI(\mul_a2/fa1_c0_r[13] ), .CO(n253), .S0(n336) );
  HS65_GS_FA1X4 U292 ( .A0(n258), .B0(n257), .CI(n256), .CO(n1648), .S0(n1644)
         );
  HS65_GS_PAOI2X1 U293 ( .A(\mul_a2/fa1_s1_r[11] ), .B(\mul_a2/fa1_s0_r[11] ), 
        .P(\mul_a2/fa1_c0_r[10] ), .Z(n259) );
  HS65_GSS_XNOR2X3 U294 ( .A(\mul_a2/fa1_c1_r[11] ), .B(n259), .Z(n322) );
  HS65_GS_IVX2 U295 ( .A(\mul_a2/fa1_c1_r[11] ), .Z(n260) );
  HS65_GS_NOR2X2 U296 ( .A(n260), .B(n259), .Z(n261) );
  HS65_GS_AOI12X2 U297 ( .A(n321), .B(n322), .C(n261), .Z(n263) );
  HS65_GS_FA1X4 U298 ( .A0(\mul_a2/fa1_s0_r[12] ), .B0(\mul_a2/fa1_s1_r[12] ), 
        .CI(\mul_a2/fa1_c0_r[11] ), .CO(n340), .S0(n321) );
  HS65_GS_FA1X4 U299 ( .A0(\mul_a2/fa1_s0_r[13] ), .B0(\mul_a2/fa1_s1_r[13] ), 
        .CI(\mul_a2/fa1_c0_r[12] ), .CO(n335), .S0(n339) );
  HS65_GSS_XOR2X3 U300 ( .A(\mul_a2/fa1_s2_r[13] ), .B(\mul_a2/fa1_c1_r[12] ), 
        .Z(n338) );
  HS65_GS_IVX2 U301 ( .A(n264), .Z(n262) );
  HS65_GS_NOR2X2 U302 ( .A(n263), .B(n262), .Z(n1119) );
  HS65_GSS_XOR2X3 U303 ( .A(n264), .B(n263), .Z(n334) );
  HS65_GSS_XOR3X2 U304 ( .A(\mul_a2/fa1_s1_r[10] ), .B(\mul_a2/fa1_c0_r[9] ), 
        .C(\mul_a2/fa1_s0_r[10] ), .Z(n304) );
  HS65_GS_PAO2X4 U305 ( .A(\mul_a2/fa1_s0_r[9] ), .B(\mul_a2/fa1_c0_r[8] ), 
        .P(\mul_a2/fa1_s1_r[9] ), .Z(n265) );
  HS65_GSS_XOR2X3 U306 ( .A(\mul_a2/fa1_c1_r[9] ), .B(n265), .Z(n305) );
  HS65_GS_NAND2X2 U307 ( .A(n304), .B(n305), .Z(n303) );
  HS65_GS_NAND2X2 U308 ( .A(\mul_a2/fa1_c1_r[9] ), .B(n265), .Z(n266) );
  HS65_GS_NAND2X2 U309 ( .A(n303), .B(n266), .Z(n271) );
  HS65_GS_IVX2 U310 ( .A(n271), .Z(n269) );
  HS65_GS_PAOI2X1 U311 ( .A(\mul_a2/fa1_s1_r[10] ), .B(\mul_a2/fa1_c0_r[9] ), 
        .P(\mul_a2/fa1_s0_r[10] ), .Z(n317) );
  HS65_GSS_XNOR2X3 U312 ( .A(\mul_a2/fa1_c1_r[10] ), .B(n317), .Z(n268) );
  HS65_GSS_XOR3X2 U313 ( .A(\mul_a2/fa1_s1_r[11] ), .B(\mul_a2/fa1_s0_r[11] ), 
        .C(\mul_a2/fa1_c0_r[10] ), .Z(n267) );
  HS65_GS_NAND2X2 U314 ( .A(n267), .B(n268), .Z(n327) );
  HS65_GS_OAI21X2 U315 ( .A(n268), .B(n267), .C(n327), .Z(n270) );
  HS65_GS_NOR2X2 U316 ( .A(n269), .B(n270), .Z(n326) );
  HS65_GSS_XOR2X3 U317 ( .A(n271), .B(n270), .Z(n316) );
  HS65_GSS_XOR3X2 U318 ( .A(\mul_a2/fa1_s1_r[8] ), .B(\mul_a2/fa1_c0_r[7] ), 
        .C(\mul_a2/fa1_s0_r[8] ), .Z(n275) );
  HS65_GS_PAO2X4 U319 ( .A(\mul_a2/fa1_s0_r[7] ), .B(\mul_a2/fa1_c0_r[6] ), 
        .P(\mul_a2/fa1_s1_r[7] ), .Z(n276) );
  HS65_GS_NAND2X2 U320 ( .A(n275), .B(n276), .Z(n274) );
  HS65_GS_PAOI2X1 U321 ( .A(\mul_a2/fa1_s1_r[8] ), .B(\mul_a2/fa1_c0_r[7] ), 
        .P(\mul_a2/fa1_s0_r[8] ), .Z(n301) );
  HS65_GSS_XNOR2X3 U322 ( .A(\mul_a2/fa1_c1_r[8] ), .B(n301), .Z(n273) );
  HS65_GSS_XOR3X2 U323 ( .A(\mul_a2/fa1_s0_r[9] ), .B(\mul_a2/fa1_c0_r[8] ), 
        .C(\mul_a2/fa1_s1_r[9] ), .Z(n272) );
  HS65_GS_NAND2X2 U324 ( .A(n272), .B(n273), .Z(n309) );
  HS65_GS_OAI21X2 U325 ( .A(n273), .B(n272), .C(n309), .Z(n300) );
  HS65_GS_NOR2X2 U326 ( .A(n274), .B(n300), .Z(n308) );
  HS65_GSS_XOR3X2 U327 ( .A(\mul_a2/fa1_s0_r[7] ), .B(\mul_a2/fa1_c0_r[6] ), 
        .C(\mul_a2/fa1_s1_r[7] ), .Z(n281) );
  HS65_GS_PAO2X4 U328 ( .A(\mul_a2/fa1_s1_r[6] ), .B(\mul_a2/fa1_s0_r[6] ), 
        .P(\mul_a2/fa1_c0_r[5] ), .Z(n282) );
  HS65_GS_NAND2X2 U329 ( .A(n281), .B(n282), .Z(n280) );
  HS65_GS_IVX2 U330 ( .A(n280), .Z(n278) );
  HS65_GS_OAI21X2 U331 ( .A(n276), .B(n275), .C(n274), .Z(n277) );
  HS65_GS_IVX2 U332 ( .A(n277), .Z(n296) );
  HS65_GS_NAND2X2 U333 ( .A(n278), .B(n296), .Z(n299) );
  HS65_GSS_XOR3X2 U334 ( .A(\mul_a2/fa1_s1_r[6] ), .B(\mul_a2/fa1_s0_r[6] ), 
        .C(\mul_a2/fa1_c0_r[5] ), .Z(n291) );
  HS65_GS_AND2X4 U335 ( .A(\mul_a2/fa1_s0_r[5] ), .B(\mul_a2/fa1_c0_r[4] ), 
        .Z(n279) );
  HS65_GS_NAND2X2 U336 ( .A(n291), .B(n279), .Z(n283) );
  HS65_GS_OAI21X2 U337 ( .A(n282), .B(n281), .C(n280), .Z(n294) );
  HS65_GS_NOR2X2 U338 ( .A(n283), .B(n294), .Z(n297) );
  HS65_GSS_XOR2X3 U339 ( .A(\mul_a2/fa1_c0_r[4] ), .B(\mul_a2/fa1_s0_r[5] ), 
        .Z(n288) );
  HS65_GS_AND2X4 U340 ( .A(\mul_a2/fa1_c0_r[3] ), .B(\mul_a2/fa1_s0_r[4] ), 
        .Z(n284) );
  HS65_GS_AND2X4 U341 ( .A(n288), .B(n284), .Z(n285) );
  HS65_GS_NAND2X2 U342 ( .A(n285), .B(n291), .Z(n293) );
  HS65_GS_AND2X4 U343 ( .A(\mul_a2/fa1_c0_r[2] ), .B(\mul_a2/fa1_s0_r[3] ), 
        .Z(n287) );
  HS65_GSS_XOR2X3 U344 ( .A(\mul_a2/fa1_c0_r[3] ), .B(\mul_a2/fa1_s0_r[4] ), 
        .Z(n286) );
  HS65_GS_AND2X4 U345 ( .A(n287), .B(n286), .Z(n289) );
  HS65_GS_AND2X4 U346 ( .A(n289), .B(n288), .Z(n290) );
  HS65_GS_NAND2X2 U347 ( .A(n291), .B(n290), .Z(n292) );
  HS65_GS_PAOI2X1 U348 ( .A(n294), .B(n293), .P(n292), .Z(n295) );
  HS65_GS_PAOI2X1 U349 ( .A(n297), .B(n296), .P(n295), .Z(n298) );
  HS65_GS_PAOI2X1 U350 ( .A(n300), .B(n299), .P(n298), .Z(n307) );
  HS65_GS_IVX2 U351 ( .A(\mul_a2/fa1_c1_r[8] ), .Z(n302) );
  HS65_GS_NOR2X2 U352 ( .A(n302), .B(n301), .Z(n312) );
  HS65_GS_OAI21X2 U353 ( .A(n305), .B(n304), .C(n303), .Z(n310) );
  HS65_GSS_XNOR2X3 U354 ( .A(n312), .B(n310), .Z(n306) );
  HS65_GS_PAOI2X1 U355 ( .A(n308), .B(n307), .P(n306), .Z(n315) );
  HS65_GS_IVX2 U356 ( .A(n309), .Z(n313) );
  HS65_GS_IVX2 U357 ( .A(n310), .Z(n311) );
  HS65_GS_OAI21X2 U358 ( .A(n313), .B(n312), .C(n311), .Z(n314) );
  HS65_GS_PAOI2X1 U359 ( .A(n316), .B(n315), .P(n314), .Z(n325) );
  HS65_GS_IVX2 U360 ( .A(\mul_a2/fa1_c1_r[10] ), .Z(n318) );
  HS65_GS_NOR2X2 U361 ( .A(n318), .B(n317), .Z(n330) );
  HS65_GS_IVX2 U362 ( .A(n330), .Z(n319) );
  HS65_GS_NAND2X2 U363 ( .A(n319), .B(n327), .Z(n323) );
  HS65_GS_NAND2X2 U364 ( .A(n321), .B(n322), .Z(n320) );
  HS65_GS_OAI21X2 U365 ( .A(n322), .B(n321), .C(n320), .Z(n328) );
  HS65_GSS_XNOR2X3 U366 ( .A(n323), .B(n328), .Z(n324) );
  HS65_GS_PAOI2X1 U367 ( .A(n326), .B(n325), .P(n324), .Z(n333) );
  HS65_GS_IVX2 U368 ( .A(n327), .Z(n331) );
  HS65_GS_IVX2 U369 ( .A(n328), .Z(n329) );
  HS65_GS_OAI21X2 U370 ( .A(n331), .B(n330), .C(n329), .Z(n332) );
  HS65_GS_PAOI2X1 U371 ( .A(n334), .B(n333), .P(n332), .Z(n1118) );
  HS65_GS_AND2X4 U372 ( .A(\mul_a2/fa1_s2_r[13] ), .B(\mul_a2/fa1_c1_r[12] ), 
        .Z(n343) );
  HS65_GS_FA1X4 U373 ( .A0(n337), .B0(n336), .CI(n335), .CO(n256), .S0(n342)
         );
  HS65_GS_FA1X4 U374 ( .A0(n340), .B0(n339), .CI(n338), .CO(n341), .S0(n264)
         );
  HS65_GS_PAO2X4 U375 ( .A(n1119), .B(n1118), .P(n1142), .Z(n1643) );
  HS65_GS_FA1X4 U376 ( .A0(n343), .B0(n342), .CI(n341), .CO(n1642), .S0(n1142)
         );
  HS65_GS_FA1X4 U377 ( .A0(n346), .B0(n345), .CI(n344), .CO(n1652), .S0(n1646)
         );
  HS65_GS_FA1X4 U378 ( .A0(n349), .B0(n348), .CI(n347), .CO(n1656), .S0(n1650)
         );
  HS65_GS_FA1X4 U379 ( .A0(n352), .B0(n351), .CI(n350), .CO(n1660), .S0(n1654)
         );
  HS65_GS_FA1X4 U380 ( .A0(n355), .B0(n354), .CI(n353), .CO(n1664), .S0(n1658)
         );
  HS65_GS_FA1X4 U381 ( .A0(n358), .B0(n357), .CI(n356), .CO(n1668), .S0(n1662)
         );
  HS65_GS_FA1X4 U382 ( .A0(n361), .B0(n360), .CI(n359), .CO(n1672), .S0(n1666)
         );
  HS65_GS_FA1X4 U383 ( .A0(n364), .B0(n363), .CI(n362), .CO(n1676), .S0(n1670)
         );
  HS65_GS_FA1X4 U384 ( .A0(\mul_a2/fa1_c1_r[21] ), .B0(\mul_a2/fa1_c2_r[21] ), 
        .CI(\mul_a2/fa1_s2_r[22] ), .CO(n373), .S0(n367) );
  HS65_GS_FA1X4 U385 ( .A0(n367), .B0(n366), .CI(n365), .CO(n372), .S0(n362)
         );
  HS65_GS_FA1X4 U386 ( .A0(n370), .B0(n369), .CI(n368), .CO(n375), .S0(n371)
         );
  HS65_GS_FA1X4 U387 ( .A0(n373), .B0(n372), .CI(n371), .CO(n1679), .S0(n1674)
         );
  HS65_GS_FA1X4 U388 ( .A0(n376), .B0(n375), .CI(n374), .CO(n1684), .S0(n1678)
         );
  HS65_GS_FA1X4 U389 ( .A0(n379), .B0(n378), .CI(n377), .CO(n1688), .S0(n1682)
         );
  HS65_GS_FA1X4 U390 ( .A0(n382), .B0(n381), .CI(n380), .CO(n1692), .S0(n1686)
         );
  HS65_GS_FA1X4 U391 ( .A0(\mul_a2/fa1_c1_r[25] ), .B0(\mul_a2/fa1_c2_r[25] ), 
        .CI(\mul_a2/fa1_s2_r[26] ), .CO(n391), .S0(n385) );
  HS65_GS_FA1X4 U392 ( .A0(n385), .B0(n384), .CI(n383), .CO(n390), .S0(n380)
         );
  HS65_GS_FA1X4 U393 ( .A0(n388), .B0(n387), .CI(n386), .CO(n393), .S0(n389)
         );
  HS65_GS_FA1X4 U394 ( .A0(n391), .B0(n390), .CI(n389), .CO(n1695), .S0(n1690)
         );
  HS65_GS_FA1X4 U395 ( .A0(n394), .B0(n393), .CI(n392), .CO(n1122), .S0(n1694)
         );
  HS65_GS_FA1X4 U396 ( .A0(n397), .B0(n396), .CI(n395), .CO(n1129), .S0(n1120)
         );
  HS65_GS_FA1X4 U397 ( .A0(n400), .B0(n399), .CI(n398), .CO(n1132), .S0(n1127)
         );
  HS65_GS_AND2X4 U398 ( .A(\mul_a2/fa1_c1_r[29] ), .B(\mul_a2/fa1_s2_r[30] ), 
        .Z(n409) );
  HS65_GS_FA1X4 U399 ( .A0(n403), .B0(n402), .CI(n401), .CO(n408), .S0(n398)
         );
  HS65_GS_FA1X4 U400 ( .A0(n406), .B0(n405), .CI(n404), .CO(n412), .S0(n407)
         );
  HS65_GS_FA1X4 U401 ( .A0(n409), .B0(n408), .CI(n407), .CO(n1124), .S0(n1130)
         );
  HS65_GS_FA1X4 U402 ( .A0(n412), .B0(n411), .CI(n410), .CO(n420), .S0(n1126)
         );
  HS65_GS_FA1X4 U403 ( .A0(n415), .B0(n414), .CI(n413), .CO(n416), .S0(n411)
         );
  HS65_GSS_XOR3X2 U404 ( .A(\mul_a2/fa1_s2_r[33] ), .B(\mul_a2/fa1_s0_r[33] ), 
        .C(n416), .Z(n418) );
  HS65_GSS_XOR2X3 U405 ( .A(\mul_a2/fa1_c1_r[32] ), .B(\mul_a2/fa1_c0_r[32] ), 
        .Z(n417) );
  HS65_GSS_XOR3X2 U406 ( .A(n418), .B(\mul_a2/fa1_s1_r[33] ), .C(n417), .Z(
        n419) );
  HS65_GSS_XOR3X2 U407 ( .A(n421), .B(n420), .C(n419), .Z(n422) );
  HS65_GSS_XOR3X2 U408 ( .A(n424), .B(n423), .C(n422), .Z(
        \mul_a2/result_sat[15] ) );
  HS65_GS_IVX2 U409 ( .A(x_z1[15]), .Z(n1492) );
  HS65_GS_AND2X4 U410 ( .A(\mul_b0/fa1_s0_r[31] ), .B(\mul_b0/fa1_s1_r[31] ), 
        .Z(n426) );
  HS65_GSS_XOR2X3 U411 ( .A(\mul_b0/fa1_s0_r[32] ), .B(\mul_b0/fa1_s1_r[32] ), 
        .Z(n425) );
  HS65_GS_AND2X4 U412 ( .A(\mul_b0/fa1_s1_r[32] ), .B(\mul_b0/fa1_s0_r[32] ), 
        .Z(n518) );
  HS65_GS_AND2X4 U413 ( .A(\mul_b0/fa1_s0_r[29] ), .B(\mul_b0/fa1_s1_r[29] ), 
        .Z(n430) );
  HS65_GSS_XOR2X3 U414 ( .A(\mul_b0/fa1_s0_r[30] ), .B(\mul_b0/fa1_s1_r[30] ), 
        .Z(n429) );
  HS65_GSS_XOR2X3 U415 ( .A(\mul_b0/fa1_s0_r[31] ), .B(\mul_b0/fa1_s1_r[31] ), 
        .Z(n428) );
  HS65_GS_AND2X4 U416 ( .A(\mul_b0/fa1_s0_r[30] ), .B(\mul_b0/fa1_s1_r[30] ), 
        .Z(n427) );
  HS65_GS_FA1X4 U417 ( .A0(\mul_b0/fa1_s2_r[32] ), .B0(n426), .CI(n425), .CO(
        n519), .S0(n515) );
  HS65_GS_FA1X4 U418 ( .A0(\mul_b0/fa1_s2_r[31] ), .B0(n428), .CI(n427), .CO(
        n514), .S0(n512) );
  HS65_GSS_XOR2X3 U419 ( .A(n515), .B(n514), .Z(n1022) );
  HS65_GS_AOI12X2 U420 ( .A(n511), .B(n512), .C(n1022), .Z(n1021) );
  HS65_GS_NAND2X2 U421 ( .A(n512), .B(n511), .Z(n510) );
  HS65_GS_IVX2 U422 ( .A(n510), .Z(n513) );
  HS65_GS_AND2X4 U423 ( .A(\mul_b0/fa1_s0_r[28] ), .B(\mul_b0/fa1_s1_r[28] ), 
        .Z(n432) );
  HS65_GSS_XOR2X3 U424 ( .A(\mul_b0/fa1_s0_r[29] ), .B(\mul_b0/fa1_s1_r[29] ), 
        .Z(n431) );
  HS65_GS_FA1X4 U425 ( .A0(\mul_b0/fa1_s2_r[30] ), .B0(n430), .CI(n429), .CO(
        n511), .S0(n1033) );
  HS65_GS_AND2X4 U426 ( .A(\mul_b0/fa1_s0_r[27] ), .B(\mul_b0/fa1_s1_r[27] ), 
        .Z(n434) );
  HS65_GSS_XOR2X3 U427 ( .A(\mul_b0/fa1_s0_r[28] ), .B(\mul_b0/fa1_s1_r[28] ), 
        .Z(n433) );
  HS65_GS_FA1X4 U428 ( .A0(\mul_b0/fa1_s2_r[29] ), .B0(n432), .CI(n431), .CO(
        n1034), .S0(n1030) );
  HS65_GS_AND2X4 U429 ( .A(\mul_b0/fa1_s0_r[26] ), .B(\mul_b0/fa1_s1_r[26] ), 
        .Z(n503) );
  HS65_GSS_XOR2X3 U430 ( .A(\mul_b0/fa1_s0_r[27] ), .B(\mul_b0/fa1_s1_r[27] ), 
        .Z(n502) );
  HS65_GS_FA1X4 U431 ( .A0(\mul_b0/fa1_s2_r[28] ), .B0(n434), .CI(n433), .CO(
        n1031), .S0(n1532) );
  HS65_GS_FA1X4 U432 ( .A0(\mul_b0/fa1_s0_r[20] ), .B0(\mul_b0/fa1_s1_r[20] ), 
        .CI(\mul_b0/fa1_c0_r[19] ), .CO(n490), .S0(n435) );
  HS65_GS_FA1X4 U433 ( .A0(\mul_b0/fa1_s0_r[19] ), .B0(\mul_b0/fa1_s1_r[19] ), 
        .CI(\mul_b0/fa1_c0_r[18] ), .CO(n436), .S0(n482) );
  HS65_GS_FA1X4 U434 ( .A0(\mul_b0/fa1_s2_r[20] ), .B0(n436), .CI(n435), .CO(
        n1549), .S0(n1552) );
  HS65_GS_FA1X4 U435 ( .A0(\mul_b0/fa1_s0_r[17] ), .B0(\mul_b0/fa1_s1_r[17] ), 
        .CI(\mul_b0/fa1_c0_r[16] ), .CO(n485), .S0(n437) );
  HS65_GS_FA1X4 U436 ( .A0(\mul_b0/fa1_s0_r[18] ), .B0(\mul_b0/fa1_s1_r[18] ), 
        .CI(\mul_b0/fa1_c0_r[17] ), .CO(n483), .S0(n484) );
  HS65_GS_FA1X4 U437 ( .A0(\mul_b0/fa1_s0_r[16] ), .B0(\mul_b0/fa1_s1_r[16] ), 
        .CI(\mul_b0/fa1_c0_r[15] ), .CO(n438), .S0(n439) );
  HS65_GS_FA1X4 U438 ( .A0(\mul_b0/fa1_s2_r[17] ), .B0(n438), .CI(n437), .CO(
        n481), .S0(n477) );
  HS65_GS_FA1X4 U439 ( .A0(\mul_b0/fa1_s0_r[15] ), .B0(\mul_b0/fa1_s1_r[15] ), 
        .CI(\mul_b0/fa1_c0_r[14] ), .CO(n440), .S0(n441) );
  HS65_GS_FA1X4 U440 ( .A0(\mul_b0/fa1_s2_r[16] ), .B0(n440), .CI(n439), .CO(
        n478), .S0(n474) );
  HS65_GS_FA1X4 U441 ( .A0(\mul_b0/fa1_s0_r[14] ), .B0(\mul_b0/fa1_s1_r[14] ), 
        .CI(\mul_b0/fa1_c0_r[13] ), .CO(n442), .S0(n443) );
  HS65_GS_FA1X4 U442 ( .A0(\mul_b0/fa1_s2_r[15] ), .B0(n442), .CI(n441), .CO(
        n475), .S0(n471) );
  HS65_GS_FA1X4 U443 ( .A0(\mul_b0/fa1_s0_r[13] ), .B0(\mul_b0/fa1_s1_r[13] ), 
        .CI(\mul_b0/fa1_c0_r[12] ), .CO(n444), .S0(n445) );
  HS65_GS_FA1X4 U444 ( .A0(\mul_b0/fa1_s2_r[14] ), .B0(n444), .CI(n443), .CO(
        n472), .S0(n468) );
  HS65_GS_FA1X4 U445 ( .A0(\mul_b0/fa1_s2_r[13] ), .B0(n446), .CI(n445), .CO(
        n469), .S0(n466) );
  HS65_GS_FA1X4 U446 ( .A0(\mul_b0/fa1_s0_r[12] ), .B0(\mul_b0/fa1_s1_r[12] ), 
        .CI(\mul_b0/fa1_c0_r[11] ), .CO(n446), .S0(n459) );
  HS65_GS_FA1X4 U447 ( .A0(\mul_b0/fa1_s0_r[11] ), .B0(\mul_b0/fa1_s1_r[11] ), 
        .CI(\mul_b0/fa1_c0_r[10] ), .CO(n458), .S0(n463) );
  HS65_GS_FA1X4 U448 ( .A0(\mul_b0/fa1_s0_r[8] ), .B0(\mul_b0/fa1_s1_r[8] ), 
        .CI(\mul_b0/fa1_c0_r[7] ), .CO(n451), .S0(n449) );
  HS65_GS_AND2X4 U449 ( .A(\mul_b0/fa1_c0_r[5] ), .B(\mul_b0/fa1_s0_r[6] ), 
        .Z(n447) );
  HS65_GS_PAO2X4 U450 ( .A(n447), .B(\mul_b0/fa1_s0_r[7] ), .P(
        \mul_b0/fa1_c0_r[6] ), .Z(n448) );
  HS65_GS_OAI112X1 U451 ( .A(n451), .B(n450), .C(n449), .D(n448), .Z(n457) );
  HS65_GS_NAND2X2 U452 ( .A(n451), .B(n450), .Z(n456) );
  HS65_GS_FA1X4 U453 ( .A0(\mul_b0/fa1_s0_r[9] ), .B0(\mul_b0/fa1_s1_r[9] ), 
        .CI(\mul_b0/fa1_c0_r[8] ), .CO(n453), .S0(n450) );
  HS65_GS_FA1X4 U454 ( .A0(\mul_b0/fa1_s0_r[10] ), .B0(\mul_b0/fa1_s1_r[10] ), 
        .CI(\mul_b0/fa1_c0_r[9] ), .CO(n462), .S0(n452) );
  HS65_GS_OAI22X1 U455 ( .A(n462), .B(n463), .C(n453), .D(n452), .Z(n455) );
  HS65_GS_OAI112X1 U456 ( .A(n462), .B(n463), .C(n453), .D(n452), .Z(n454) );
  HS65_GS_CBI4I1X3 U457 ( .A(n457), .B(n456), .C(n455), .D(n454), .Z(n461) );
  HS65_GS_FA1X4 U458 ( .A0(\mul_b0/fa1_s2_r[12] ), .B0(n459), .CI(n458), .CO(
        n465), .S0(n460) );
  HS65_GS_CB4I1X4 U459 ( .A(n463), .B(n462), .C(n461), .D(n460), .Z(n464) );
  HS65_GS_PAOI2X1 U460 ( .A(n466), .B(n465), .P(n464), .Z(n1070) );
  HS65_GS_NAND2X2 U461 ( .A(n468), .B(n469), .Z(n467) );
  HS65_GS_OAI21X2 U462 ( .A(n468), .B(n469), .C(n467), .Z(n1069) );
  HS65_GS_NOR2X2 U463 ( .A(n1070), .B(n1069), .Z(n1068) );
  HS65_GS_AOI12X2 U464 ( .A(n469), .B(n468), .C(n1068), .Z(n1066) );
  HS65_GS_NAND2X2 U465 ( .A(n471), .B(n472), .Z(n470) );
  HS65_GS_OAI21X2 U466 ( .A(n471), .B(n472), .C(n470), .Z(n1065) );
  HS65_GS_NOR2X2 U467 ( .A(n1066), .B(n1065), .Z(n1064) );
  HS65_GS_AOI12X2 U468 ( .A(n472), .B(n471), .C(n1064), .Z(n1062) );
  HS65_GS_NAND2X2 U469 ( .A(n474), .B(n475), .Z(n473) );
  HS65_GS_OAI21X2 U470 ( .A(n474), .B(n475), .C(n473), .Z(n1061) );
  HS65_GS_NOR2X2 U471 ( .A(n1062), .B(n1061), .Z(n1060) );
  HS65_GS_AOI12X2 U472 ( .A(n475), .B(n474), .C(n1060), .Z(n1058) );
  HS65_GS_NAND2X2 U473 ( .A(n477), .B(n478), .Z(n476) );
  HS65_GS_OAI21X2 U474 ( .A(n477), .B(n478), .C(n476), .Z(n1057) );
  HS65_GS_NOR2X2 U475 ( .A(n1058), .B(n1057), .Z(n1056) );
  HS65_GS_AOI12X2 U476 ( .A(n478), .B(n477), .C(n1056), .Z(n1054) );
  HS65_GS_NAND2X2 U477 ( .A(n480), .B(n481), .Z(n479) );
  HS65_GS_OAI21X2 U478 ( .A(n480), .B(n481), .C(n479), .Z(n1053) );
  HS65_GS_NOR2X2 U479 ( .A(n1054), .B(n1053), .Z(n1052) );
  HS65_GS_AOI12X2 U480 ( .A(n481), .B(n480), .C(n1052), .Z(n1559) );
  HS65_GS_FA1X4 U481 ( .A0(\mul_b0/fa1_s2_r[19] ), .B0(n483), .CI(n482), .CO(
        n1553), .S0(n487) );
  HS65_GS_FA1X4 U482 ( .A0(\mul_b0/fa1_s2_r[18] ), .B0(n485), .CI(n484), .CO(
        n486), .S0(n480) );
  HS65_GS_NAND2X2 U483 ( .A(n487), .B(n486), .Z(n488) );
  HS65_GS_OAI21X2 U484 ( .A(n487), .B(n486), .C(n488), .Z(n1560) );
  HS65_GS_OAI21X2 U485 ( .A(n1559), .B(n1560), .C(n488), .Z(n1551) );
  HS65_GS_FA1X4 U486 ( .A0(\mul_b0/fa1_s2_r[21] ), .B0(n490), .CI(n489), .CO(
        n1544), .S0(n1548) );
  HS65_GS_FA1X4 U487 ( .A0(\mul_b0/fa1_s0_r[21] ), .B0(\mul_b0/fa1_s1_r[21] ), 
        .CI(\mul_b0/fa1_c0_r[20] ), .CO(n492), .S0(n489) );
  HS65_GSS_XOR2X3 U488 ( .A(\mul_b0/fa1_s0_r[22] ), .B(\mul_b0/fa1_s1_r[22] ), 
        .Z(n491) );
  HS65_GS_FA1X4 U489 ( .A0(\mul_b0/fa1_s2_r[22] ), .B0(n492), .CI(n491), .CO(
        n1540), .S0(n1543) );
  HS65_GS_AND2X4 U490 ( .A(\mul_b0/fa1_s1_r[22] ), .B(\mul_b0/fa1_s0_r[22] ), 
        .Z(n494) );
  HS65_GSS_XOR2X3 U491 ( .A(\mul_b0/fa1_s0_r[23] ), .B(\mul_b0/fa1_s1_r[23] ), 
        .Z(n493) );
  HS65_GS_FA1X4 U492 ( .A0(\mul_b0/fa1_s2_r[23] ), .B0(n494), .CI(n493), .CO(
        n1536), .S0(n1539) );
  HS65_GS_AND2X4 U493 ( .A(\mul_b0/fa1_s1_r[23] ), .B(\mul_b0/fa1_s0_r[23] ), 
        .Z(n496) );
  HS65_GSS_XOR2X3 U494 ( .A(\mul_b0/fa1_s0_r[24] ), .B(\mul_b0/fa1_s1_r[24] ), 
        .Z(n495) );
  HS65_GS_AND2X4 U495 ( .A(\mul_b0/fa1_s1_r[24] ), .B(\mul_b0/fa1_s0_r[24] ), 
        .Z(n498) );
  HS65_GSS_XOR2X3 U496 ( .A(\mul_b0/fa1_s0_r[25] ), .B(\mul_b0/fa1_s1_r[25] ), 
        .Z(n497) );
  HS65_GS_FA1X4 U497 ( .A0(\mul_b0/fa1_s2_r[24] ), .B0(n496), .CI(n495), .CO(
        n1047), .S0(n1535) );
  HS65_GS_PAOI2X1 U498 ( .A(n1050), .B(n1048), .P(n1047), .Z(n1045) );
  HS65_GS_AND2X4 U499 ( .A(\mul_b0/fa1_s1_r[25] ), .B(\mul_b0/fa1_s0_r[25] ), 
        .Z(n505) );
  HS65_GSS_XOR2X3 U500 ( .A(\mul_b0/fa1_s0_r[26] ), .B(\mul_b0/fa1_s1_r[26] ), 
        .Z(n504) );
  HS65_GS_FA1X4 U501 ( .A0(\mul_b0/fa1_s2_r[25] ), .B0(n498), .CI(n497), .CO(
        n499), .S0(n1048) );
  HS65_GS_NAND2X2 U502 ( .A(n500), .B(n499), .Z(n501) );
  HS65_GS_OAI21X2 U503 ( .A(n500), .B(n499), .C(n501), .Z(n1046) );
  HS65_GS_OA12X4 U504 ( .A(n1045), .B(n1046), .C(n501), .Z(n1042) );
  HS65_GS_FA1X4 U505 ( .A0(\mul_b0/fa1_s2_r[27] ), .B0(n503), .CI(n502), .CO(
        n1533), .S0(n507) );
  HS65_GS_FA1X4 U506 ( .A0(\mul_b0/fa1_s2_r[26] ), .B0(n505), .CI(n504), .CO(
        n506), .S0(n500) );
  HS65_GS_NAND2X2 U507 ( .A(n507), .B(n506), .Z(n508) );
  HS65_GS_OAI21X2 U508 ( .A(n507), .B(n506), .C(n508), .Z(n1043) );
  HS65_GS_OAI21X2 U509 ( .A(n1042), .B(n1043), .C(n508), .Z(n1531) );
  HS65_GS_IVX2 U510 ( .A(n509), .Z(n1028) );
  HS65_GS_OAI21X2 U511 ( .A(n512), .B(n511), .C(n510), .Z(n1027) );
  HS65_GS_NOR2X2 U512 ( .A(n1028), .B(n1027), .Z(n1026) );
  HS65_GS_AOI12X2 U513 ( .A(n1022), .B(n513), .C(n1026), .Z(n1025) );
  HS65_GS_NAND2X2 U514 ( .A(n515), .B(n514), .Z(n516) );
  HS65_GS_OAI21X2 U515 ( .A(n1021), .B(n1025), .C(n516), .Z(n517) );
  HS65_GSS_XOR3X2 U516 ( .A(n519), .B(n518), .C(n517), .Z(n520) );
  HS65_GSS_XOR2X3 U517 ( .A(\mul_b0/fa1_s2_r[33] ), .B(n520), .Z(n521) );
  HS65_GSS_XOR3X2 U518 ( .A(\mul_b0/fa1_s0_r[33] ), .B(\mul_b0/fa1_s1_r[33] ), 
        .C(n521), .Z(\mul_b0/result_sat[15] ) );
  HS65_GS_BFX4 U519 ( .A(valid_in), .Z(n1406) );
  HS65_GS_BFX4 U520 ( .A(n1406), .Z(n1892) );
  HS65_GS_AND2X4 U521 ( .A(\mul_a1/fa1_s0_r[32] ), .B(\mul_a1/fa1_s1_r[32] ), 
        .Z(n744) );
  HS65_GSS_XOR2X3 U522 ( .A(\mul_a1/fa1_s1_r[31] ), .B(\mul_a1/fa1_s0_r[31] ), 
        .Z(n731) );
  HS65_GS_AND2X4 U523 ( .A(\mul_a1/fa1_s0_r[30] ), .B(\mul_a1/fa1_s1_r[30] ), 
        .Z(n730) );
  HS65_GSS_XOR2X3 U524 ( .A(\mul_a1/fa1_s1_r[32] ), .B(\mul_a1/fa1_s0_r[32] ), 
        .Z(n523) );
  HS65_GS_AND2X4 U525 ( .A(\mul_a1/fa1_s0_r[31] ), .B(\mul_a1/fa1_s1_r[31] ), 
        .Z(n522) );
  HS65_GS_AND2X4 U526 ( .A(n736), .B(n735), .Z(n525) );
  HS65_GS_FA1X4 U527 ( .A0(n523), .B0(\mul_a1/fa1_s2_r[32] ), .CI(n522), .CO(
        n524), .S0(n735) );
  HS65_GSS_XOR2X3 U528 ( .A(n525), .B(n524), .Z(n741) );
  HS65_GSS_XOR2X3 U529 ( .A(\mul_a1/fa1_s1_r[29] ), .B(\mul_a1/fa1_s0_r[29] ), 
        .Z(n533) );
  HS65_GS_AND2X4 U530 ( .A(\mul_a1/fa1_s0_r[28] ), .B(\mul_a1/fa1_s1_r[28] ), 
        .Z(n532) );
  HS65_GSS_XOR2X3 U531 ( .A(\mul_a1/fa1_s2_r[29] ), .B(\mul_a1/fa1_c2_r[28] ), 
        .Z(n531) );
  HS65_GS_AOI12X2 U532 ( .A(\mul_a1/fa1_c2_r[28] ), .B(\mul_a1/fa1_s2_r[29] ), 
        .C(n528), .Z(n529) );
  HS65_GS_AND2X4 U533 ( .A(\mul_a1/fa1_s0_r[29] ), .B(\mul_a1/fa1_s1_r[29] ), 
        .Z(n734) );
  HS65_GSS_XOR2X3 U534 ( .A(\mul_a1/fa1_s1_r[30] ), .B(\mul_a1/fa1_s0_r[30] ), 
        .Z(n733) );
  HS65_GSS_XOR2X3 U535 ( .A(\mul_a1/fa1_s2_r[30] ), .B(\mul_a1/fa1_c2_r[29] ), 
        .Z(n732) );
  HS65_GS_AND2X4 U536 ( .A(\mul_a1/fa1_s2_r[29] ), .B(\mul_a1/fa1_c2_r[28] ), 
        .Z(n527) );
  HS65_GS_NAND3X2 U537 ( .A(n533), .B(n532), .C(n527), .Z(n526) );
  HS65_GS_OAI21X2 U538 ( .A(n528), .B(n527), .C(n526), .Z(n728) );
  HS65_GS_NOR2X2 U539 ( .A(n729), .B(n728), .Z(n727) );
  HS65_GS_NOR2X2 U540 ( .A(n529), .B(n727), .Z(n1079) );
  HS65_GSS_XOR2X3 U541 ( .A(\mul_a1/fa1_s1_r[28] ), .B(\mul_a1/fa1_s0_r[28] ), 
        .Z(n542) );
  HS65_GS_AND2X4 U542 ( .A(\mul_a1/fa1_s0_r[27] ), .B(\mul_a1/fa1_s1_r[27] ), 
        .Z(n530) );
  HS65_GS_FA1X4 U543 ( .A0(\mul_a1/fa1_c2_r[27] ), .B0(\mul_a1/fa1_s2_r[28] ), 
        .CI(n530), .CO(n536), .S0(n543) );
  HS65_GS_AOI12X2 U544 ( .A(n542), .B(n543), .C(n536), .Z(n537) );
  HS65_GS_FA1X4 U545 ( .A0(n533), .B0(n532), .CI(n531), .CO(n528), .S0(n726)
         );
  HS65_GS_NAND2X2 U546 ( .A(n543), .B(n542), .Z(n541) );
  HS65_GS_IVX2 U547 ( .A(n541), .Z(n535) );
  HS65_GS_NAND3X2 U548 ( .A(\mul_a1/fa1_c2_r[27] ), .B(\mul_a1/fa1_s2_r[28] ), 
        .C(n535), .Z(n534) );
  HS65_GS_OAI21X2 U549 ( .A(n536), .B(n535), .C(n534), .Z(n725) );
  HS65_GS_NOR2X2 U550 ( .A(n726), .B(n725), .Z(n724) );
  HS65_GS_NOR2X2 U551 ( .A(n537), .B(n724), .Z(n1085) );
  HS65_GS_AND2X4 U552 ( .A(\mul_a1/fa1_s1_r[26] ), .B(\mul_a1/fa1_s0_r[26] ), 
        .Z(n538) );
  HS65_GSS_XOR2X3 U553 ( .A(\mul_a1/fa1_s1_r[27] ), .B(\mul_a1/fa1_s0_r[27] ), 
        .Z(n715) );
  HS65_GS_NAND2X2 U554 ( .A(n716), .B(n715), .Z(n714) );
  HS65_GS_IVX2 U555 ( .A(n714), .Z(n540) );
  HS65_GS_FA1X4 U556 ( .A0(\mul_a1/fa1_c2_r[26] ), .B0(\mul_a1/fa1_s2_r[27] ), 
        .CI(n538), .CO(n539), .S0(n716) );
  HS65_GS_AOI12X2 U557 ( .A(n715), .B(n716), .C(n539), .Z(n544) );
  HS65_GS_AOI13X2 U558 ( .A(n540), .B(\mul_a1/fa1_c2_r[26] ), .C(
        \mul_a1/fa1_s2_r[27] ), .D(n544), .Z(n723) );
  HS65_GS_OAI21X2 U559 ( .A(n543), .B(n542), .C(n541), .Z(n722) );
  HS65_GS_NAND2X2 U560 ( .A(n723), .B(n722), .Z(n721) );
  HS65_GS_NOR2AX3 U561 ( .A(n721), .B(n544), .Z(n1075) );
  HS65_GS_AND2X4 U562 ( .A(\mul_a1/fa1_s1_r[24] ), .B(\mul_a1/fa1_s0_r[24] ), 
        .Z(n545) );
  HS65_GSS_XOR2X3 U563 ( .A(\mul_a1/fa1_s1_r[25] ), .B(\mul_a1/fa1_s0_r[25] ), 
        .Z(n553) );
  HS65_GS_NAND2X2 U564 ( .A(n554), .B(n553), .Z(n552) );
  HS65_GS_IVX2 U565 ( .A(n552), .Z(n547) );
  HS65_GS_FA1X4 U566 ( .A0(\mul_a1/fa1_c2_r[24] ), .B0(\mul_a1/fa1_s2_r[25] ), 
        .CI(n545), .CO(n546), .S0(n554) );
  HS65_GS_NOR2X2 U567 ( .A(n547), .B(n546), .Z(n548) );
  HS65_GS_AOI13X2 U568 ( .A(n547), .B(\mul_a1/fa1_c2_r[24] ), .C(
        \mul_a1/fa1_s2_r[25] ), .D(n548), .Z(n707) );
  HS65_GS_AND2X4 U569 ( .A(\mul_a1/fa1_s0_r[25] ), .B(\mul_a1/fa1_s1_r[25] ), 
        .Z(n709) );
  HS65_GSS_XOR2X3 U570 ( .A(\mul_a1/fa1_s0_r[26] ), .B(\mul_a1/fa1_s1_r[26] ), 
        .Z(n712) );
  HS65_GS_NAND2X2 U571 ( .A(n711), .B(n712), .Z(n708) );
  HS65_GS_OAI21X2 U572 ( .A(n711), .B(n712), .C(n708), .Z(n706) );
  HS65_GS_NAND2X2 U573 ( .A(n707), .B(n706), .Z(n705) );
  HS65_GS_NOR2AX3 U574 ( .A(n705), .B(n548), .Z(n1574) );
  HS65_GS_AND2X4 U575 ( .A(\mul_a1/fa1_s1_r[23] ), .B(\mul_a1/fa1_s0_r[23] ), 
        .Z(n549) );
  HS65_GSS_XOR2X3 U576 ( .A(\mul_a1/fa1_s0_r[24] ), .B(\mul_a1/fa1_s1_r[24] ), 
        .Z(n696) );
  HS65_GS_NAND2X2 U577 ( .A(n697), .B(n696), .Z(n695) );
  HS65_GS_IVX2 U578 ( .A(n695), .Z(n551) );
  HS65_GS_FA1X4 U579 ( .A0(\mul_a1/fa1_c2_r[23] ), .B0(\mul_a1/fa1_s2_r[24] ), 
        .CI(n549), .CO(n550), .S0(n697) );
  HS65_GS_AOI12X2 U580 ( .A(n696), .B(n697), .C(n550), .Z(n555) );
  HS65_GS_AOI13X2 U581 ( .A(n551), .B(\mul_a1/fa1_s2_r[24] ), .C(
        \mul_a1/fa1_c2_r[23] ), .D(n555), .Z(n557) );
  HS65_GS_OAI21X2 U582 ( .A(n554), .B(n553), .C(n552), .Z(n556) );
  HS65_GS_AOI12X2 U583 ( .A(n557), .B(n556), .C(n555), .Z(n1570) );
  HS65_GSS_XNOR2X3 U584 ( .A(n557), .B(n556), .Z(n1117) );
  HS65_GS_IVX2 U585 ( .A(n1117), .Z(n704) );
  HS65_GSS_XOR2X3 U586 ( .A(\mul_a1/fa1_s1_r[22] ), .B(\mul_a1/fa1_s0_r[22] ), 
        .Z(n567) );
  HS65_GS_PAO2X4 U587 ( .A(\mul_a1/fa1_s1_r[21] ), .B(\mul_a1/fa1_s0_r[21] ), 
        .P(\mul_a1/fa1_c0_r[20] ), .Z(n558) );
  HS65_GS_FA1X4 U588 ( .A0(\mul_a1/fa1_c2_r[21] ), .B0(\mul_a1/fa1_s2_r[22] ), 
        .CI(n558), .CO(n559), .S0(n568) );
  HS65_GS_AOI12X2 U589 ( .A(n567), .B(n568), .C(n559), .Z(n562) );
  HS65_GS_NAND2X2 U590 ( .A(n568), .B(n567), .Z(n566) );
  HS65_GS_IVX2 U591 ( .A(n566), .Z(n560) );
  HS65_GS_AOI13X2 U592 ( .A(n560), .B(\mul_a1/fa1_s2_r[22] ), .C(
        \mul_a1/fa1_c2_r[21] ), .D(n562), .Z(n686) );
  HS65_GS_AND2X4 U593 ( .A(\mul_a1/fa1_s0_r[22] ), .B(\mul_a1/fa1_s1_r[22] ), 
        .Z(n691) );
  HS65_GSS_XOR2X3 U594 ( .A(\mul_a1/fa1_s0_r[23] ), .B(\mul_a1/fa1_s1_r[23] ), 
        .Z(n693) );
  HS65_GS_NAND2X2 U595 ( .A(n692), .B(n693), .Z(n690) );
  HS65_GS_OAI21X2 U596 ( .A(n692), .B(n693), .C(n690), .Z(n685) );
  HS65_GS_AND2X4 U597 ( .A(n686), .B(n685), .Z(n561) );
  HS65_GS_NOR2X2 U598 ( .A(n562), .B(n561), .Z(n688) );
  HS65_GSS_XOR3X2 U599 ( .A(\mul_a1/fa1_s1_r[21] ), .B(\mul_a1/fa1_s0_r[21] ), 
        .C(\mul_a1/fa1_c0_r[20] ), .Z(n581) );
  HS65_GS_PAO2X4 U600 ( .A(\mul_a1/fa1_s1_r[20] ), .B(\mul_a1/fa1_s0_r[20] ), 
        .P(\mul_a1/fa1_c0_r[19] ), .Z(n563) );
  HS65_GS_FA1X4 U601 ( .A0(\mul_a1/fa1_c2_r[20] ), .B0(\mul_a1/fa1_s2_r[21] ), 
        .CI(n563), .CO(n564), .S0(n582) );
  HS65_GS_AOI12X2 U602 ( .A(n581), .B(n582), .C(n564), .Z(n570) );
  HS65_GS_NAND2X2 U603 ( .A(n582), .B(n581), .Z(n580) );
  HS65_GS_IVX2 U604 ( .A(n580), .Z(n565) );
  HS65_GS_AOI13X2 U605 ( .A(n565), .B(\mul_a1/fa1_s2_r[21] ), .C(
        \mul_a1/fa1_c2_r[20] ), .D(n570), .Z(n679) );
  HS65_GS_OAI21X2 U606 ( .A(n568), .B(n567), .C(n566), .Z(n678) );
  HS65_GS_AND2X4 U607 ( .A(n679), .B(n678), .Z(n569) );
  HS65_GS_NOR2X2 U608 ( .A(n570), .B(n569), .Z(n684) );
  HS65_GS_PAO2X4 U609 ( .A(\mul_a1/fa1_s1_r[18] ), .B(\mul_a1/fa1_s0_r[18] ), 
        .P(\mul_a1/fa1_c0_r[17] ), .Z(n571) );
  HS65_GSS_XOR3X2 U610 ( .A(\mul_a1/fa1_c0_r[18] ), .B(\mul_a1/fa1_s1_r[19] ), 
        .C(\mul_a1/fa1_s0_r[19] ), .Z(n589) );
  HS65_GS_NAND2X2 U611 ( .A(n590), .B(n589), .Z(n588) );
  HS65_GS_IVX2 U612 ( .A(n588), .Z(n574) );
  HS65_GS_FA1X4 U613 ( .A0(\mul_a1/fa1_c2_r[18] ), .B0(\mul_a1/fa1_s2_r[19] ), 
        .CI(n571), .CO(n573), .S0(n590) );
  HS65_GS_NOR2X2 U614 ( .A(n574), .B(n573), .Z(n572) );
  HS65_GS_AOI13X2 U615 ( .A(n574), .B(\mul_a1/fa1_c2_r[18] ), .C(
        \mul_a1/fa1_s2_r[19] ), .D(n572), .Z(n677) );
  HS65_GS_PAO2X4 U616 ( .A(\mul_a1/fa1_c0_r[18] ), .B(\mul_a1/fa1_s1_r[19] ), 
        .P(\mul_a1/fa1_s0_r[19] ), .Z(n576) );
  HS65_GSS_XOR3X2 U617 ( .A(\mul_a1/fa1_s1_r[20] ), .B(\mul_a1/fa1_s0_r[20] ), 
        .C(\mul_a1/fa1_c0_r[19] ), .Z(n578) );
  HS65_GS_NAND2X2 U618 ( .A(n577), .B(n578), .Z(n575) );
  HS65_GS_OAI21X2 U619 ( .A(n577), .B(n578), .C(n575), .Z(n676) );
  HS65_GS_NAND2X2 U620 ( .A(n677), .B(n676), .Z(n675) );
  HS65_GS_OAI21X2 U621 ( .A(n574), .B(n573), .C(n675), .Z(n1858) );
  HS65_GS_IVX2 U622 ( .A(n575), .Z(n682) );
  HS65_GS_FA1X4 U623 ( .A0(\mul_a1/fa1_c2_r[19] ), .B0(\mul_a1/fa1_s2_r[20] ), 
        .CI(n576), .CO(n681), .S0(n577) );
  HS65_GS_AOI12X2 U624 ( .A(n578), .B(n577), .C(n681), .Z(n579) );
  HS65_GS_AOI13X2 U625 ( .A(n682), .B(\mul_a1/fa1_s2_r[20] ), .C(
        \mul_a1/fa1_c2_r[19] ), .D(n579), .Z(n584) );
  HS65_GS_OAI21X2 U626 ( .A(n582), .B(n581), .C(n580), .Z(n583) );
  HS65_GS_NAND2X2 U627 ( .A(n584), .B(n583), .Z(n680) );
  HS65_GS_OA12X4 U628 ( .A(n584), .B(n583), .C(n680), .Z(n1857) );
  HS65_GS_PAO2X4 U629 ( .A(\mul_a1/fa1_s1_r[17] ), .B(\mul_a1/fa1_s0_r[17] ), 
        .P(\mul_a1/fa1_c0_r[16] ), .Z(n585) );
  HS65_GSS_XOR3X2 U630 ( .A(\mul_a1/fa1_s1_r[18] ), .B(\mul_a1/fa1_s0_r[18] ), 
        .C(\mul_a1/fa1_c0_r[17] ), .Z(n660) );
  HS65_GS_NAND2X2 U631 ( .A(n661), .B(n660), .Z(n659) );
  HS65_GS_IVX2 U632 ( .A(n659), .Z(n587) );
  HS65_GS_FA1X4 U633 ( .A0(\mul_a1/fa1_c2_r[17] ), .B0(\mul_a1/fa1_s2_r[18] ), 
        .CI(n585), .CO(n586), .S0(n661) );
  HS65_GS_AOI12X2 U634 ( .A(n660), .B(n661), .C(n586), .Z(n591) );
  HS65_GS_AOI13X2 U635 ( .A(n587), .B(\mul_a1/fa1_s2_r[18] ), .C(
        \mul_a1/fa1_c2_r[17] ), .D(n591), .Z(n673) );
  HS65_GS_OAI21X2 U636 ( .A(n590), .B(n589), .C(n588), .Z(n672) );
  HS65_GS_AO12X4 U637 ( .A(n673), .B(n672), .C(n591), .Z(n1854) );
  HS65_GS_PAO2X4 U638 ( .A(\mul_a1/fa1_s1_r[14] ), .B(\mul_a1/fa1_s0_r[14] ), 
        .P(\mul_a1/fa1_c0_r[13] ), .Z(n638) );
  HS65_GS_NAND2X2 U639 ( .A(\mul_a1/fa1_s2_r[15] ), .B(\mul_a1/fa1_c2_r[14] ), 
        .Z(n636) );
  HS65_GS_OAI21X2 U640 ( .A(\mul_a1/fa1_s2_r[15] ), .B(\mul_a1/fa1_c2_r[14] ), 
        .C(n636), .Z(n592) );
  HS65_GSS_XOR3X2 U641 ( .A(\mul_a1/fa1_c0_r[14] ), .B(\mul_a1/fa1_s1_r[15] ), 
        .C(\mul_a1/fa1_s0_r[15] ), .Z(n640) );
  HS65_GS_NAND2AX4 U642 ( .A(n592), .B(n640), .Z(n634) );
  HS65_GS_NAND2AX4 U643 ( .A(n640), .B(n592), .Z(n633) );
  HS65_GS_NAND2X2 U644 ( .A(n634), .B(n633), .Z(n593) );
  HS65_GSS_XNOR2X3 U645 ( .A(n638), .B(n593), .Z(n594) );
  HS65_GSS_XOR3X2 U646 ( .A(\mul_a1/fa1_s1_r[14] ), .B(\mul_a1/fa1_s0_r[14] ), 
        .C(\mul_a1/fa1_c0_r[13] ), .Z(n597) );
  HS65_GS_PAO2X4 U647 ( .A(\mul_a1/fa1_c0_r[12] ), .B(\mul_a1/fa1_s1_r[13] ), 
        .P(\mul_a1/fa1_s0_r[13] ), .Z(n596) );
  HS65_GS_AND2X4 U648 ( .A(n594), .B(n595), .Z(n1566) );
  HS65_GSS_XOR2X3 U649 ( .A(n595), .B(n594), .Z(n1562) );
  HS65_GS_PAO2X4 U650 ( .A(\mul_a1/fa1_c0_r[11] ), .B(\mul_a1/fa1_s1_r[12] ), 
        .P(\mul_a1/fa1_s0_r[12] ), .Z(n599) );
  HS65_GSS_XOR3X2 U651 ( .A(\mul_a1/fa1_c0_r[12] ), .B(\mul_a1/fa1_s1_r[13] ), 
        .C(\mul_a1/fa1_s0_r[13] ), .Z(n598) );
  HS65_GS_FA1X4 U652 ( .A0(\mul_a1/fa1_s2_r[14] ), .B0(n597), .CI(n596), .CO(
        n595), .S0(n631) );
  HS65_GS_FA1X4 U653 ( .A0(\mul_a1/fa1_s2_r[13] ), .B0(n599), .CI(n598), .CO(
        n632), .S0(n628) );
  HS65_GSS_XNOR3X2 U654 ( .A(\mul_a1/fa1_c0_r[11] ), .B(\mul_a1/fa1_s1_r[12] ), 
        .C(\mul_a1/fa1_s0_r[12] ), .Z(n600) );
  HS65_GS_PAOI2X1 U655 ( .A(\mul_a1/fa1_s1_r[11] ), .B(\mul_a1/fa1_c0_r[10] ), 
        .P(\mul_a1/fa1_s0_r[11] ), .Z(n601) );
  HS65_GS_NOR2X2 U656 ( .A(n600), .B(n601), .Z(n627) );
  HS65_GSS_XNOR3X2 U657 ( .A(\mul_a1/fa1_s1_r[11] ), .B(\mul_a1/fa1_c0_r[10] ), 
        .C(\mul_a1/fa1_s0_r[11] ), .Z(n602) );
  HS65_GS_PAOI2X1 U658 ( .A(\mul_a1/fa1_s1_r[10] ), .B(\mul_a1/fa1_c0_r[9] ), 
        .P(\mul_a1/fa1_s0_r[10] ), .Z(n603) );
  HS65_GS_NOR2X2 U659 ( .A(n602), .B(n603), .Z(n625) );
  HS65_GSS_XOR2X3 U660 ( .A(n601), .B(n600), .Z(n624) );
  HS65_GSS_XNOR3X2 U661 ( .A(\mul_a1/fa1_s1_r[10] ), .B(\mul_a1/fa1_c0_r[9] ), 
        .C(\mul_a1/fa1_s0_r[10] ), .Z(n604) );
  HS65_GS_PAOI2X1 U662 ( .A(\mul_a1/fa1_s1_r[9] ), .B(\mul_a1/fa1_c0_r[8] ), 
        .P(\mul_a1/fa1_s0_r[9] ), .Z(n605) );
  HS65_GS_NOR2X2 U663 ( .A(n604), .B(n605), .Z(n622) );
  HS65_GSS_XOR2X3 U664 ( .A(n603), .B(n602), .Z(n621) );
  HS65_GSS_XNOR3X2 U665 ( .A(\mul_a1/fa1_s1_r[9] ), .B(\mul_a1/fa1_c0_r[8] ), 
        .C(\mul_a1/fa1_s0_r[9] ), .Z(n606) );
  HS65_GS_PAOI2X1 U666 ( .A(\mul_a1/fa1_s1_r[8] ), .B(\mul_a1/fa1_c0_r[7] ), 
        .P(\mul_a1/fa1_s0_r[8] ), .Z(n607) );
  HS65_GS_NOR2X2 U667 ( .A(n606), .B(n607), .Z(n619) );
  HS65_GSS_XOR2X3 U668 ( .A(n605), .B(n604), .Z(n618) );
  HS65_GSS_XOR2X3 U669 ( .A(n607), .B(n606), .Z(n616) );
  HS65_GSS_XNOR3X2 U670 ( .A(\mul_a1/fa1_s1_r[8] ), .B(\mul_a1/fa1_c0_r[7] ), 
        .C(\mul_a1/fa1_s0_r[8] ), .Z(n611) );
  HS65_GS_NAND2X2 U671 ( .A(\mul_a1/fa1_c0_r[6] ), .B(\mul_a1/fa1_s0_r[7] ), 
        .Z(n608) );
  HS65_GS_NOR2X2 U672 ( .A(n611), .B(n608), .Z(n615) );
  HS65_GSS_XNOR2X3 U673 ( .A(\mul_a1/fa1_c0_r[6] ), .B(\mul_a1/fa1_s0_r[7] ), 
        .Z(n610) );
  HS65_GS_NAND2X2 U674 ( .A(\mul_a1/fa1_c0_r[5] ), .B(\mul_a1/fa1_s0_r[6] ), 
        .Z(n609) );
  HS65_GS_NOR2X2 U675 ( .A(n610), .B(n609), .Z(n613) );
  HS65_GS_IVX2 U676 ( .A(n611), .Z(n612) );
  HS65_GS_AND2X4 U677 ( .A(n613), .B(n612), .Z(n614) );
  HS65_GS_PAO2X4 U678 ( .A(n616), .B(n615), .P(n614), .Z(n617) );
  HS65_GS_PAO2X4 U679 ( .A(n619), .B(n618), .P(n617), .Z(n620) );
  HS65_GS_PAO2X4 U680 ( .A(n622), .B(n621), .P(n620), .Z(n623) );
  HS65_GS_PAO2X4 U681 ( .A(n625), .B(n624), .P(n623), .Z(n626) );
  HS65_GS_PAOI2X1 U682 ( .A(n628), .B(n627), .P(n626), .Z(n1094) );
  HS65_GS_NAND2X2 U683 ( .A(n631), .B(n632), .Z(n629) );
  HS65_GS_OAI21X2 U684 ( .A(n631), .B(n632), .C(n629), .Z(n1093) );
  HS65_GS_NOR2X2 U685 ( .A(n1094), .B(n1093), .Z(n630) );
  HS65_GS_AO12X4 U686 ( .A(n632), .B(n631), .C(n630), .Z(n1561) );
  HS65_GS_AND2X4 U687 ( .A(n1562), .B(n1561), .Z(n1565) );
  HS65_GS_IVX2 U688 ( .A(n636), .Z(n639) );
  HS65_GS_NAND2X2 U689 ( .A(n638), .B(n633), .Z(n635) );
  HS65_GS_NAND3X2 U690 ( .A(n636), .B(n635), .C(n634), .Z(n644) );
  HS65_GS_IVX2 U691 ( .A(n644), .Z(n637) );
  HS65_GS_AOI13X2 U692 ( .A(n640), .B(n639), .C(n638), .D(n637), .Z(n642) );
  HS65_GS_PAO2X4 U693 ( .A(\mul_a1/fa1_c0_r[14] ), .B(\mul_a1/fa1_s1_r[15] ), 
        .P(\mul_a1/fa1_s0_r[15] ), .Z(n646) );
  HS65_GSS_XOR3X2 U694 ( .A(\mul_a1/fa1_c0_r[15] ), .B(\mul_a1/fa1_s1_r[16] ), 
        .C(\mul_a1/fa1_s0_r[16] ), .Z(n648) );
  HS65_GS_NAND2X2 U695 ( .A(n647), .B(n648), .Z(n645) );
  HS65_GS_OAI21X2 U696 ( .A(n647), .B(n648), .C(n645), .Z(n641) );
  HS65_GS_NAND2X2 U697 ( .A(n642), .B(n641), .Z(n643) );
  HS65_GS_OAI21X2 U698 ( .A(n642), .B(n641), .C(n643), .Z(n1564) );
  HS65_GS_NAND2X2 U699 ( .A(n644), .B(n643), .Z(n650) );
  HS65_GS_NOR2AX3 U700 ( .A(n651), .B(n650), .Z(n653) );
  HS65_GS_IVX2 U701 ( .A(n645), .Z(n666) );
  HS65_GS_FA1X4 U702 ( .A0(\mul_a1/fa1_c2_r[15] ), .B0(\mul_a1/fa1_s2_r[16] ), 
        .CI(n646), .CO(n665), .S0(n647) );
  HS65_GS_AOI12X2 U703 ( .A(n648), .B(n647), .C(n665), .Z(n649) );
  HS65_GS_AOI13X2 U704 ( .A(n666), .B(\mul_a1/fa1_s2_r[16] ), .C(
        \mul_a1/fa1_c2_r[15] ), .D(n649), .Z(n663) );
  HS65_GS_PAO2X4 U705 ( .A(\mul_a1/fa1_c0_r[15] ), .B(\mul_a1/fa1_s1_r[16] ), 
        .P(\mul_a1/fa1_s0_r[16] ), .Z(n655) );
  HS65_GSS_XOR3X2 U706 ( .A(\mul_a1/fa1_s1_r[17] ), .B(\mul_a1/fa1_s0_r[17] ), 
        .C(\mul_a1/fa1_c0_r[16] ), .Z(n657) );
  HS65_GS_NAND2X2 U707 ( .A(n656), .B(n657), .Z(n654) );
  HS65_GS_OAI21X2 U708 ( .A(n656), .B(n657), .C(n654), .Z(n662) );
  HS65_GSS_XOR2X3 U709 ( .A(n663), .B(n662), .Z(n1096) );
  HS65_GSS_XOR2X3 U710 ( .A(n651), .B(n650), .Z(n1097) );
  HS65_GS_NOR2X2 U711 ( .A(n1096), .B(n1097), .Z(n652) );
  HS65_GS_NOR2X2 U712 ( .A(n653), .B(n652), .Z(n1099) );
  HS65_GS_IVX2 U713 ( .A(n654), .Z(n671) );
  HS65_GS_FA1X4 U714 ( .A0(\mul_a1/fa1_c2_r[16] ), .B0(\mul_a1/fa1_s2_r[17] ), 
        .CI(n655), .CO(n670), .S0(n656) );
  HS65_GS_AOI12X2 U715 ( .A(n657), .B(n656), .C(n670), .Z(n658) );
  HS65_GS_AOI13X2 U716 ( .A(n671), .B(\mul_a1/fa1_s2_r[17] ), .C(
        \mul_a1/fa1_c2_r[16] ), .D(n658), .Z(n668) );
  HS65_GS_OAI21X2 U717 ( .A(n661), .B(n660), .C(n659), .Z(n667) );
  HS65_GSS_XOR2X3 U718 ( .A(n668), .B(n667), .Z(n1101) );
  HS65_GS_NAND2X2 U719 ( .A(n663), .B(n662), .Z(n664) );
  HS65_GS_OAI21X2 U720 ( .A(n666), .B(n665), .C(n664), .Z(n1098) );
  HS65_GS_PAOI2X1 U721 ( .A(n1099), .B(n1101), .P(n1098), .Z(n1104) );
  HS65_GS_NAND2X2 U722 ( .A(n668), .B(n667), .Z(n669) );
  HS65_GS_OA12X4 U723 ( .A(n671), .B(n670), .C(n669), .Z(n1103) );
  HS65_GSS_XOR2X3 U724 ( .A(n673), .B(n672), .Z(n1106) );
  HS65_GS_IVX2 U725 ( .A(n1106), .Z(n674) );
  HS65_GS_PAOI2X1 U726 ( .A(n1104), .B(n1103), .P(n674), .Z(n1853) );
  HS65_GS_OA12X4 U727 ( .A(n677), .B(n676), .C(n675), .Z(n1852) );
  HS65_GSS_XOR2X3 U728 ( .A(n679), .B(n678), .Z(n1111) );
  HS65_GS_OAI21X2 U729 ( .A(n682), .B(n681), .C(n680), .Z(n1108) );
  HS65_GS_PAOI2X1 U730 ( .A(n1109), .B(n1111), .P(n1108), .Z(n683) );
  HS65_GS_NOR2X2 U731 ( .A(n684), .B(n683), .Z(n687) );
  HS65_GSS_XNOR2X3 U732 ( .A(n684), .B(n683), .Z(n1862) );
  HS65_GSS_XNOR2X3 U733 ( .A(n686), .B(n685), .Z(n1861) );
  HS65_GS_NOR2X2 U734 ( .A(n1862), .B(n1861), .Z(n1860) );
  HS65_GS_NOR2X2 U735 ( .A(n687), .B(n1860), .Z(n689) );
  HS65_GS_NOR2X2 U736 ( .A(n688), .B(n689), .Z(n698) );
  HS65_GSS_XNOR2X3 U737 ( .A(n689), .B(n688), .Z(n1866) );
  HS65_GS_IVX2 U738 ( .A(n690), .Z(n703) );
  HS65_GS_FA1X4 U739 ( .A0(\mul_a1/fa1_c2_r[22] ), .B0(\mul_a1/fa1_s2_r[23] ), 
        .CI(n691), .CO(n702), .S0(n692) );
  HS65_GS_AOI12X2 U740 ( .A(n693), .B(n692), .C(n702), .Z(n694) );
  HS65_GS_AOI13X2 U741 ( .A(n703), .B(\mul_a1/fa1_s2_r[23] ), .C(
        \mul_a1/fa1_c2_r[22] ), .D(n694), .Z(n700) );
  HS65_GS_OAI21X2 U742 ( .A(n697), .B(n696), .C(n695), .Z(n699) );
  HS65_GSS_XNOR2X3 U743 ( .A(n700), .B(n699), .Z(n1865) );
  HS65_GS_NOR2X2 U744 ( .A(n1866), .B(n1865), .Z(n1864) );
  HS65_GS_OR2X4 U745 ( .A(n698), .B(n1864), .Z(n1114) );
  HS65_GS_NAND2X2 U746 ( .A(n700), .B(n699), .Z(n701) );
  HS65_GS_OAI21X2 U747 ( .A(n703), .B(n702), .C(n701), .Z(n1113) );
  HS65_GS_PAOI2X1 U748 ( .A(n704), .B(n1114), .P(n1113), .Z(n1569) );
  HS65_GS_OAI21X2 U749 ( .A(n707), .B(n706), .C(n705), .Z(n1568) );
  HS65_GS_IVX2 U750 ( .A(n708), .Z(n713) );
  HS65_GS_FA1X4 U751 ( .A0(\mul_a1/fa1_c2_r[25] ), .B0(\mul_a1/fa1_s2_r[26] ), 
        .CI(n709), .CO(n710), .S0(n711) );
  HS65_GS_AOI12X2 U752 ( .A(n712), .B(n711), .C(n710), .Z(n719) );
  HS65_GS_AOI13X2 U753 ( .A(n713), .B(\mul_a1/fa1_c2_r[25] ), .C(
        \mul_a1/fa1_s2_r[26] ), .D(n719), .Z(n718) );
  HS65_GS_OAI21X2 U754 ( .A(n716), .B(n715), .C(n714), .Z(n717) );
  HS65_GS_NAND2X2 U755 ( .A(n718), .B(n717), .Z(n720) );
  HS65_GS_OAI21X2 U756 ( .A(n718), .B(n717), .C(n720), .Z(n1572) );
  HS65_GS_NOR2AX3 U757 ( .A(n720), .B(n719), .Z(n1577) );
  HS65_GS_OAI21X2 U758 ( .A(n723), .B(n722), .C(n721), .Z(n1576) );
  HS65_GS_AO12X4 U759 ( .A(n726), .B(n725), .C(n724), .Z(n1073) );
  HS65_GS_AO12X4 U760 ( .A(n729), .B(n728), .C(n727), .Z(n1083) );
  HS65_GS_AND2X4 U761 ( .A(\mul_a1/fa1_s2_r[30] ), .B(\mul_a1/fa1_c2_r[29] ), 
        .Z(n739) );
  HS65_GS_FA1X4 U762 ( .A0(\mul_a1/fa1_s2_r[31] ), .B0(n731), .CI(n730), .CO(
        n736), .S0(n738) );
  HS65_GS_FA1X4 U763 ( .A0(n734), .B0(n733), .CI(n732), .CO(n737), .S0(n729)
         );
  HS65_GSS_XOR2X3 U764 ( .A(n736), .B(n735), .Z(n1081) );
  HS65_GS_FA1X4 U765 ( .A0(n739), .B0(n738), .CI(n737), .CO(n1080), .S0(n1077)
         );
  HS65_GSS_XOR2X3 U766 ( .A(n741), .B(n740), .Z(n742) );
  HS65_GSS_XOR3X2 U767 ( .A(n742), .B(\mul_a1/fa1_s0_r[33] ), .C(
        \mul_a1/fa1_s1_r[33] ), .Z(n743) );
  HS65_GSS_XOR3X2 U768 ( .A(n744), .B(\mul_a1/fa1_s2_r[33] ), .C(n743), .Z(
        \mul_a1/result_sat[15] ) );
  HS65_GS_IVX4 U769 ( .A(y_z1[15]), .Z(n1815) );
  HS65_GS_IVX2 U770 ( .A(y_z1[14]), .Z(n1817) );
  HS65_GS_IVX2 U771 ( .A(y_z1[13]), .Z(n1819) );
  HS65_GS_IVX2 U772 ( .A(y_z1[12]), .Z(n1821) );
  HS65_GS_IVX2 U773 ( .A(y_z1[11]), .Z(n1823) );
  HS65_GS_IVX2 U774 ( .A(y_z1[10]), .Z(n1825) );
  HS65_GS_IVX2 U775 ( .A(y_z1[9]), .Z(n1827) );
  HS65_GS_IVX2 U776 ( .A(y_z1[8]), .Z(n1829) );
  HS65_GS_IVX2 U777 ( .A(y_z1[7]), .Z(n1831) );
  HS65_GS_IVX2 U778 ( .A(y_z1[6]), .Z(n1833) );
  HS65_GS_IVX2 U779 ( .A(y_z1[5]), .Z(n1835) );
  HS65_GS_IVX2 U780 ( .A(y_z1[4]), .Z(n1837) );
  HS65_GS_IVX2 U781 ( .A(y_z1[3]), .Z(n1839) );
  HS65_GS_IVX2 U782 ( .A(y_z1[2]), .Z(n1841) );
  HS65_GS_IVX2 U783 ( .A(y_z1[1]), .Z(n1843) );
  HS65_GS_IVX2 U784 ( .A(y_z1[0]), .Z(n1842) );
  HS65_GS_NOR2X2 U785 ( .A(y_z1[15]), .B(n1813), .Z(n1886) );
  HS65_GS_FA1X4 U786 ( .A0(\mul_b2/fa1_s0_r[32] ), .B0(\mul_b2/fa1_s1_r[32] ), 
        .CI(\mul_b2/fa1_c0_r[31] ), .CO(n863), .S0(n745) );
  HS65_GS_FA1X4 U787 ( .A0(\mul_b2/fa1_s0_r[31] ), .B0(\mul_b2/fa1_s1_r[31] ), 
        .CI(\mul_b2/fa1_c0_r[30] ), .CO(n746), .S0(n748) );
  HS65_GS_FA1X4 U788 ( .A0(\mul_b2/fa1_s0_r[30] ), .B0(\mul_b2/fa1_s1_r[30] ), 
        .CI(\mul_b2/fa1_c0_r[29] ), .CO(n747), .S0(n749) );
  HS65_GS_FA1X4 U789 ( .A0(\mul_b2/fa1_s2_r[32] ), .B0(n746), .CI(n745), .CO(
        n864), .S0(n860) );
  HS65_GS_FA1X4 U790 ( .A0(\mul_b2/fa1_s2_r[31] ), .B0(n748), .CI(n747), .CO(
        n859), .S0(n857) );
  HS65_GSS_XOR2X3 U791 ( .A(n860), .B(n859), .Z(n1144) );
  HS65_GS_AOI12X2 U792 ( .A(n856), .B(n857), .C(n1144), .Z(n1143) );
  HS65_GS_NAND2X2 U793 ( .A(n857), .B(n856), .Z(n855) );
  HS65_GS_IVX2 U794 ( .A(n855), .Z(n858) );
  HS65_GS_FA1X4 U795 ( .A0(\mul_b2/fa1_s0_r[29] ), .B0(\mul_b2/fa1_s1_r[29] ), 
        .CI(\mul_b2/fa1_c0_r[28] ), .CO(n750), .S0(n751) );
  HS65_GS_FA1X4 U796 ( .A0(\mul_b2/fa1_s2_r[30] ), .B0(n750), .CI(n749), .CO(
        n856), .S0(n1155) );
  HS65_GS_FA1X4 U797 ( .A0(\mul_b2/fa1_s0_r[28] ), .B0(\mul_b2/fa1_s1_r[28] ), 
        .CI(\mul_b2/fa1_c0_r[27] ), .CO(n752), .S0(n753) );
  HS65_GS_FA1X4 U798 ( .A0(\mul_b2/fa1_s2_r[29] ), .B0(n752), .CI(n751), .CO(
        n1156), .S0(n1152) );
  HS65_GS_FA1X4 U799 ( .A0(\mul_b2/fa1_s0_r[27] ), .B0(\mul_b2/fa1_s1_r[27] ), 
        .CI(\mul_b2/fa1_c0_r[26] ), .CO(n754), .S0(n847) );
  HS65_GS_FA1X4 U800 ( .A0(\mul_b2/fa1_s2_r[28] ), .B0(n754), .CI(n753), .CO(
        n1153), .S0(n1804) );
  HS65_GS_FA1X4 U801 ( .A0(\mul_b2/fa1_s0_r[25] ), .B0(\mul_b2/fa1_s1_r[25] ), 
        .CI(\mul_b2/fa1_c0_r[24] ), .CO(n850), .S0(n755) );
  HS65_GS_FA1X4 U802 ( .A0(\mul_b2/fa1_s0_r[26] ), .B0(\mul_b2/fa1_s1_r[26] ), 
        .CI(\mul_b2/fa1_c0_r[25] ), .CO(n848), .S0(n849) );
  HS65_GS_FA1X4 U803 ( .A0(\mul_b2/fa1_s0_r[24] ), .B0(\mul_b2/fa1_s1_r[24] ), 
        .CI(\mul_b2/fa1_c0_r[23] ), .CO(n756), .S0(n757) );
  HS65_GS_FA1X4 U804 ( .A0(\mul_b2/fa1_s2_r[25] ), .B0(n756), .CI(n755), .CO(
        n846), .S0(n842) );
  HS65_GS_FA1X4 U805 ( .A0(\mul_b2/fa1_s0_r[23] ), .B0(\mul_b2/fa1_s1_r[23] ), 
        .CI(\mul_b2/fa1_c0_r[22] ), .CO(n758), .S0(n759) );
  HS65_GS_FA1X4 U806 ( .A0(\mul_b2/fa1_s2_r[24] ), .B0(n758), .CI(n757), .CO(
        n843), .S0(n839) );
  HS65_GS_FA1X4 U807 ( .A0(\mul_b2/fa1_s0_r[22] ), .B0(\mul_b2/fa1_s1_r[22] ), 
        .CI(\mul_b2/fa1_c0_r[21] ), .CO(n760), .S0(n761) );
  HS65_GS_FA1X4 U808 ( .A0(\mul_b2/fa1_s2_r[23] ), .B0(n760), .CI(n759), .CO(
        n840), .S0(n836) );
  HS65_GS_FA1X4 U809 ( .A0(\mul_b2/fa1_s0_r[21] ), .B0(\mul_b2/fa1_s1_r[21] ), 
        .CI(\mul_b2/fa1_c0_r[20] ), .CO(n762), .S0(n763) );
  HS65_GS_FA1X4 U810 ( .A0(\mul_b2/fa1_s2_r[22] ), .B0(n762), .CI(n761), .CO(
        n837), .S0(n833) );
  HS65_GS_FA1X4 U811 ( .A0(\mul_b2/fa1_s0_r[20] ), .B0(\mul_b2/fa1_s1_r[20] ), 
        .CI(\mul_b2/fa1_c0_r[19] ), .CO(n764), .S0(n765) );
  HS65_GS_FA1X4 U812 ( .A0(\mul_b2/fa1_s2_r[21] ), .B0(n764), .CI(n763), .CO(
        n834), .S0(n830) );
  HS65_GS_FA1X4 U813 ( .A0(\mul_b2/fa1_s0_r[19] ), .B0(\mul_b2/fa1_s1_r[19] ), 
        .CI(\mul_b2/fa1_c0_r[18] ), .CO(n766), .S0(n768) );
  HS65_GS_FA1X4 U814 ( .A0(\mul_b2/fa1_s2_r[20] ), .B0(n766), .CI(n765), .CO(
        n831), .S0(n827) );
  HS65_GS_FA1X4 U815 ( .A0(\mul_b2/fa1_s0_r[18] ), .B0(\mul_b2/fa1_s1_r[18] ), 
        .CI(\mul_b2/fa1_c0_r[17] ), .CO(n767), .S0(n769) );
  HS65_GS_FA1X4 U816 ( .A0(\mul_b2/fa1_s2_r[19] ), .B0(n768), .CI(n767), .CO(
        n828), .S0(n824) );
  HS65_GS_FA1X4 U817 ( .A0(\mul_b2/fa1_s0_r[17] ), .B0(\mul_b2/fa1_s1_r[17] ), 
        .CI(\mul_b2/fa1_c0_r[16] ), .CO(n770), .S0(n772) );
  HS65_GS_FA1X4 U818 ( .A0(\mul_b2/fa1_s2_r[18] ), .B0(n770), .CI(n769), .CO(
        n825), .S0(n821) );
  HS65_GS_NOR2X2 U819 ( .A(n822), .B(n821), .Z(n771) );
  HS65_GS_AOI12X2 U820 ( .A(n821), .B(n822), .C(n771), .Z(n1179) );
  HS65_GS_FA1X4 U821 ( .A0(\mul_b2/fa1_s0_r[16] ), .B0(\mul_b2/fa1_s1_r[16] ), 
        .CI(\mul_b2/fa1_c0_r[15] ), .CO(n773), .S0(n775) );
  HS65_GS_FA1X4 U822 ( .A0(\mul_b2/fa1_s2_r[17] ), .B0(n773), .CI(n772), .CO(
        n822), .S0(n818) );
  HS65_GS_FA1X4 U823 ( .A0(\mul_b2/fa1_s0_r[15] ), .B0(\mul_b2/fa1_s1_r[15] ), 
        .CI(\mul_b2/fa1_c0_r[14] ), .CO(n774), .S0(n777) );
  HS65_GS_FA1X4 U824 ( .A0(\mul_b2/fa1_s2_r[16] ), .B0(n775), .CI(n774), .CO(
        n819), .S0(n815) );
  HS65_GS_NOR2X2 U825 ( .A(n816), .B(n815), .Z(n776) );
  HS65_GS_AOI12X2 U826 ( .A(n815), .B(n816), .C(n776), .Z(n1172) );
  HS65_GS_FA1X4 U827 ( .A0(\mul_b2/fa1_s0_r[14] ), .B0(\mul_b2/fa1_s1_r[14] ), 
        .CI(\mul_b2/fa1_c0_r[13] ), .CO(n778), .S0(n780) );
  HS65_GS_FA1X4 U828 ( .A0(\mul_b2/fa1_s2_r[15] ), .B0(n778), .CI(n777), .CO(
        n816), .S0(n812) );
  HS65_GS_NOR2X2 U829 ( .A(n813), .B(n812), .Z(n779) );
  HS65_GS_AOI12X2 U830 ( .A(n812), .B(n813), .C(n779), .Z(n1169) );
  HS65_GS_FA1X4 U831 ( .A0(\mul_b2/fa1_s0_r[13] ), .B0(\mul_b2/fa1_s1_r[13] ), 
        .CI(\mul_b2/fa1_c0_r[12] ), .CO(n781), .S0(n782) );
  HS65_GS_FA1X4 U832 ( .A0(\mul_b2/fa1_s2_r[14] ), .B0(n781), .CI(n780), .CO(
        n813), .S0(n809) );
  HS65_GS_FA1X4 U833 ( .A0(\mul_b2/fa1_s2_r[13] ), .B0(n783), .CI(n782), .CO(
        n810), .S0(n807) );
  HS65_GS_FA1X4 U834 ( .A0(\mul_b2/fa1_s0_r[12] ), .B0(\mul_b2/fa1_s1_r[12] ), 
        .CI(\mul_b2/fa1_c0_r[11] ), .CO(n783), .S0(n784) );
  HS65_GS_FA1X4 U835 ( .A0(\mul_b2/fa1_s2_r[12] ), .B0(n785), .CI(n784), .CO(
        n806), .S0(n804) );
  HS65_GS_FA1X4 U836 ( .A0(\mul_b2/fa1_s0_r[11] ), .B0(\mul_b2/fa1_s1_r[11] ), 
        .CI(\mul_b2/fa1_c0_r[10] ), .CO(n785), .S0(n802) );
  HS65_GS_OR2X4 U837 ( .A(\mul_b2/fa1_c0_r[6] ), .B(\mul_b2/fa1_s0_r[7] ), .Z(
        n791) );
  HS65_GS_OAI22X1 U838 ( .A(\mul_b2/fa1_c0_r[6] ), .B(\mul_b2/fa1_s0_r[7] ), 
        .C(\mul_b2/fa1_c0_r[5] ), .D(\mul_b2/fa1_s0_r[6] ), .Z(n789) );
  HS65_GS_AND2X4 U839 ( .A(\mul_b2/fa1_s0_r[3] ), .B(\mul_b2/fa1_c0_r[2] ), 
        .Z(n786) );
  HS65_GS_PAO2X4 U840 ( .A(\mul_b2/fa1_s0_r[4] ), .B(\mul_b2/fa1_c0_r[3] ), 
        .P(n786), .Z(n787) );
  HS65_GS_PAOI2X1 U841 ( .A(\mul_b2/fa1_s0_r[5] ), .B(n787), .P(
        \mul_b2/fa1_c0_r[4] ), .Z(n788) );
  HS65_GS_NOR2X2 U842 ( .A(n789), .B(n788), .Z(n790) );
  HS65_GS_AO31X4 U843 ( .A(\mul_b2/fa1_c0_r[5] ), .B(\mul_b2/fa1_s0_r[6] ), 
        .C(n791), .D(n790), .Z(n793) );
  HS65_GS_FA1X4 U844 ( .A0(\mul_b2/fa1_s0_r[8] ), .B0(\mul_b2/fa1_s1_r[8] ), 
        .CI(\mul_b2/fa1_c0_r[7] ), .CO(n795), .S0(n792) );
  HS65_GS_CB4I1X4 U845 ( .A(\mul_b2/fa1_s0_r[7] ), .B(\mul_b2/fa1_c0_r[6] ), 
        .C(n793), .D(n792), .Z(n794) );
  HS65_GS_PAO2X4 U846 ( .A(n796), .B(n795), .P(n794), .Z(n799) );
  HS65_GS_FA1X4 U847 ( .A0(\mul_b2/fa1_s0_r[10] ), .B0(\mul_b2/fa1_s1_r[10] ), 
        .CI(\mul_b2/fa1_c0_r[9] ), .CO(n801), .S0(n798) );
  HS65_GS_FA1X4 U848 ( .A0(\mul_b2/fa1_s0_r[9] ), .B0(\mul_b2/fa1_s1_r[9] ), 
        .CI(\mul_b2/fa1_c0_r[8] ), .CO(n797), .S0(n796) );
  HS65_GS_PAO2X4 U849 ( .A(n799), .B(n798), .P(n797), .Z(n800) );
  HS65_GS_PAOI2X1 U850 ( .A(n802), .B(n801), .P(n800), .Z(n803) );
  HS65_GS_NOR2AX3 U851 ( .A(n804), .B(n803), .Z(n805) );
  HS65_GS_PAOI2X1 U852 ( .A(n807), .B(n806), .P(n805), .Z(n1165) );
  HS65_GS_NAND2X2 U853 ( .A(n809), .B(n810), .Z(n808) );
  HS65_GS_OAI21X2 U854 ( .A(n809), .B(n810), .C(n808), .Z(n1164) );
  HS65_GS_NOR2X2 U855 ( .A(n1165), .B(n1164), .Z(n1163) );
  HS65_GS_AOI12X2 U856 ( .A(n810), .B(n809), .C(n1163), .Z(n1168) );
  HS65_GS_NAND2X2 U857 ( .A(n1169), .B(n1168), .Z(n811) );
  HS65_GS_OAI21X2 U858 ( .A(n813), .B(n812), .C(n811), .Z(n1171) );
  HS65_GS_NAND2X2 U859 ( .A(n1172), .B(n1171), .Z(n814) );
  HS65_GS_OAI21X2 U860 ( .A(n816), .B(n815), .C(n814), .Z(n1175) );
  HS65_GS_NAND2X2 U861 ( .A(n818), .B(n819), .Z(n817) );
  HS65_GS_OAI21X2 U862 ( .A(n818), .B(n819), .C(n817), .Z(n1174) );
  HS65_GS_NOR2X2 U863 ( .A(n1175), .B(n1174), .Z(n1173) );
  HS65_GS_AOI12X2 U864 ( .A(n819), .B(n818), .C(n1173), .Z(n1178) );
  HS65_GS_NAND2X2 U865 ( .A(n1179), .B(n1178), .Z(n820) );
  HS65_GS_OAI21X2 U866 ( .A(n822), .B(n821), .C(n820), .Z(n1182) );
  HS65_GS_NAND2X2 U867 ( .A(n824), .B(n825), .Z(n823) );
  HS65_GS_OAI21X2 U868 ( .A(n824), .B(n825), .C(n823), .Z(n1181) );
  HS65_GS_NOR2X2 U869 ( .A(n1182), .B(n1181), .Z(n1180) );
  HS65_GS_AOI12X2 U870 ( .A(n825), .B(n824), .C(n1180), .Z(n1186) );
  HS65_GS_NAND2X2 U871 ( .A(n827), .B(n828), .Z(n826) );
  HS65_GS_OAI21X2 U872 ( .A(n827), .B(n828), .C(n826), .Z(n1185) );
  HS65_GS_NOR2X2 U873 ( .A(n1186), .B(n1185), .Z(n1184) );
  HS65_GS_AOI12X2 U874 ( .A(n828), .B(n827), .C(n1184), .Z(n1190) );
  HS65_GS_NAND2X2 U875 ( .A(n830), .B(n831), .Z(n829) );
  HS65_GS_OAI21X2 U876 ( .A(n830), .B(n831), .C(n829), .Z(n1189) );
  HS65_GS_NOR2X2 U877 ( .A(n1190), .B(n1189), .Z(n1188) );
  HS65_GS_AOI12X2 U878 ( .A(n831), .B(n830), .C(n1188), .Z(n1194) );
  HS65_GS_NAND2X2 U879 ( .A(n833), .B(n834), .Z(n832) );
  HS65_GS_OAI21X2 U880 ( .A(n833), .B(n834), .C(n832), .Z(n1193) );
  HS65_GS_NOR2X2 U881 ( .A(n1194), .B(n1193), .Z(n1192) );
  HS65_GS_AOI12X2 U882 ( .A(n834), .B(n833), .C(n1192), .Z(n1198) );
  HS65_GS_NAND2X2 U883 ( .A(n836), .B(n837), .Z(n835) );
  HS65_GS_OAI21X2 U884 ( .A(n836), .B(n837), .C(n835), .Z(n1197) );
  HS65_GS_NOR2X2 U885 ( .A(n1198), .B(n1197), .Z(n1196) );
  HS65_GS_AOI12X2 U886 ( .A(n837), .B(n836), .C(n1196), .Z(n1202) );
  HS65_GS_NAND2X2 U887 ( .A(n839), .B(n840), .Z(n838) );
  HS65_GS_OAI21X2 U888 ( .A(n839), .B(n840), .C(n838), .Z(n1201) );
  HS65_GS_NOR2X2 U889 ( .A(n1202), .B(n1201), .Z(n1200) );
  HS65_GS_AOI12X2 U890 ( .A(n840), .B(n839), .C(n1200), .Z(n1206) );
  HS65_GS_NAND2X2 U891 ( .A(n842), .B(n843), .Z(n841) );
  HS65_GS_OAI21X2 U892 ( .A(n842), .B(n843), .C(n841), .Z(n1205) );
  HS65_GS_NOR2X2 U893 ( .A(n1206), .B(n1205), .Z(n1204) );
  HS65_GS_AOI12X2 U894 ( .A(n843), .B(n842), .C(n1204), .Z(n1210) );
  HS65_GS_NAND2X2 U895 ( .A(n845), .B(n846), .Z(n844) );
  HS65_GS_OAI21X2 U896 ( .A(n845), .B(n846), .C(n844), .Z(n1209) );
  HS65_GS_NOR2X2 U897 ( .A(n1210), .B(n1209), .Z(n1208) );
  HS65_GS_AOI12X2 U898 ( .A(n846), .B(n845), .C(n1208), .Z(n1801) );
  HS65_GS_FA1X4 U899 ( .A0(\mul_b2/fa1_s2_r[27] ), .B0(n848), .CI(n847), .CO(
        n1805), .S0(n852) );
  HS65_GS_FA1X4 U900 ( .A0(\mul_b2/fa1_s2_r[26] ), .B0(n850), .CI(n849), .CO(
        n851), .S0(n845) );
  HS65_GS_NAND2X2 U901 ( .A(n852), .B(n851), .Z(n853) );
  HS65_GS_OAI21X2 U902 ( .A(n852), .B(n851), .C(n853), .Z(n1802) );
  HS65_GS_OAI21X2 U903 ( .A(n1801), .B(n1802), .C(n853), .Z(n1803) );
  HS65_GS_IVX2 U904 ( .A(n854), .Z(n1150) );
  HS65_GS_OAI21X2 U905 ( .A(n857), .B(n856), .C(n855), .Z(n1149) );
  HS65_GS_NOR2X2 U906 ( .A(n1150), .B(n1149), .Z(n1148) );
  HS65_GS_AOI12X2 U907 ( .A(n1144), .B(n858), .C(n1148), .Z(n1147) );
  HS65_GS_NAND2X2 U908 ( .A(n860), .B(n859), .Z(n861) );
  HS65_GS_OAI21X2 U909 ( .A(n1143), .B(n1147), .C(n861), .Z(n862) );
  HS65_GSS_XOR3X2 U910 ( .A(n864), .B(n863), .C(n862), .Z(n865) );
  HS65_GSS_XOR3X2 U911 ( .A(\mul_b2/fa1_c0_r[32] ), .B(\mul_b2/fa1_s2_r[33] ), 
        .C(n865), .Z(n866) );
  HS65_GSS_XOR3X2 U912 ( .A(\mul_b2/fa1_s0_r[33] ), .B(\mul_b2/fa1_s1_r[33] ), 
        .C(n866), .Z(\mul_b2/result_sat[15] ) );
  HS65_GS_IVX2 U913 ( .A(x_z2[15]), .Z(n1810) );
  HS65_GS_IVX2 U914 ( .A(x_reg2[15]), .Z(n1409) );
  HS65_GS_IVX4 U915 ( .A(n1409), .Z(n1889) );
  HS65_GS_IVX2 U916 ( .A(x_reg2[1]), .Z(n1846) );
  HS65_GS_IVX2 U917 ( .A(x_reg2[3]), .Z(n1845) );
  HS65_GS_NOR2X2 U918 ( .A(n1846), .B(n1845), .Z(\mul_b2/fa1_c0[3] ) );
  HS65_GS_AOI12X2 U919 ( .A(n1846), .B(n1845), .C(\mul_b2/fa1_c0[3] ), .Z(
        \mul_b2/fa1_s0[3] ) );
  HS65_GS_IVX2 U920 ( .A(y_z2[15]), .Z(n1398) );
  HS65_GS_IVX2 U921 ( .A(y_z2[14]), .Z(n1726) );
  HS65_GS_IVX2 U922 ( .A(y_z2[13]), .Z(n1724) );
  HS65_GS_IVX2 U923 ( .A(y_z2[12]), .Z(n1722) );
  HS65_GS_IVX2 U924 ( .A(y_z2[11]), .Z(n1720) );
  HS65_GS_IVX2 U925 ( .A(y_z2[10]), .Z(n1718) );
  HS65_GS_IVX2 U926 ( .A(y_z2[9]), .Z(n1716) );
  HS65_GS_IVX2 U927 ( .A(y_z2[8]), .Z(n1714) );
  HS65_GS_IVX2 U928 ( .A(y_z2[7]), .Z(n1712) );
  HS65_GS_IVX2 U929 ( .A(y_z2[6]), .Z(n1710) );
  HS65_GS_IVX2 U930 ( .A(y_z2[5]), .Z(n1708) );
  HS65_GS_IVX2 U931 ( .A(y_z2[4]), .Z(n1706) );
  HS65_GS_IVX2 U932 ( .A(y_z2[3]), .Z(n1704) );
  HS65_GS_IVX2 U933 ( .A(y_z2[2]), .Z(n1702) );
  HS65_GS_IVX2 U934 ( .A(\mul_a2/fa1_s0[1] ), .Z(n1844) );
  HS65_GS_IVX2 U935 ( .A(\mul_a2/fa1_s0[0] ), .Z(n1314) );
  HS65_GS_IVX2 U936 ( .A(n867), .Z(n920) );
  HS65_GS_AND2X4 U937 ( .A(p_b1[1]), .B(p_b0[1]), .Z(n915) );
  HS65_GSS_XOR2X3 U938 ( .A(p_b1[1]), .B(p_b0[1]), .Z(n918) );
  HS65_GS_FA1X4 U939 ( .A0(p_b2[0]), .B0(p_b0[0]), .CI(p_b1[0]), .CO(n917), 
        .S0(n867) );
  HS65_GS_FA1X4 U940 ( .A0(p_b0[2]), .B0(p_b1[2]), .CI(p_b2[2]), .CO(n911), 
        .S0(n913) );
  HS65_GS_FA1X4 U941 ( .A0(p_b0[3]), .B0(p_b1[3]), .CI(p_b2[3]), .CO(n907), 
        .S0(n909) );
  HS65_GS_FA1X4 U942 ( .A0(p_b0[4]), .B0(p_b1[4]), .CI(p_b2[4]), .CO(n903), 
        .S0(n905) );
  HS65_GS_FA1X4 U943 ( .A0(p_b0[5]), .B0(p_b1[5]), .CI(p_b2[5]), .CO(n899), 
        .S0(n901) );
  HS65_GS_FA1X4 U944 ( .A0(p_b0[6]), .B0(p_b1[6]), .CI(p_b2[6]), .CO(n895), 
        .S0(n897) );
  HS65_GS_FA1X4 U945 ( .A0(p_b0[7]), .B0(p_b1[7]), .CI(p_b2[7]), .CO(n891), 
        .S0(n893) );
  HS65_GS_FA1X4 U946 ( .A0(p_b0[8]), .B0(p_b1[8]), .CI(p_b2[8]), .CO(n887), 
        .S0(n889) );
  HS65_GS_FA1X4 U947 ( .A0(p_b0[9]), .B0(p_b1[9]), .CI(p_b2[9]), .CO(n883), 
        .S0(n885) );
  HS65_GS_FA1X4 U948 ( .A0(p_b0[10]), .B0(p_b1[10]), .CI(p_b2[10]), .CO(n875), 
        .S0(n881) );
  HS65_GS_FA1X4 U949 ( .A0(p_b0[11]), .B0(p_b1[11]), .CI(p_b2[11]), .CO(n879), 
        .S0(n873) );
  HS65_GS_FA1X4 U950 ( .A0(p_b0[12]), .B0(p_b1[12]), .CI(p_b2[12]), .CO(n871), 
        .S0(n877) );
  HS65_GS_FA1X4 U951 ( .A0(p_b0[13]), .B0(p_b1[13]), .CI(p_b2[13]), .CO(n968), 
        .S0(n869) );
  HS65_GS_FA1X4 U952 ( .A0(p_b0[14]), .B0(p_b1[14]), .CI(p_b2[14]), .CO(n975), 
        .S0(n966) );
  HS65_GS_IVX2 U953 ( .A(p_b0[15]), .Z(n976) );
  HS65_GS_NAND2X2 U954 ( .A(p_b2[15]), .B(p_b1[15]), .Z(n977) );
  HS65_GS_OAI21X2 U955 ( .A(p_b2[15]), .B(p_b1[15]), .C(n977), .Z(n868) );
  HS65_GS_MUXI21X2 U956 ( .D0(p_b0[15]), .D1(n976), .S0(n868), .Z(n973) );
  HS65_GS_FA1X4 U957 ( .A0(n871), .B0(n870), .CI(n869), .CO(n967), .S0(n872)
         );
  HS65_GS_IVX2 U958 ( .A(n872), .Z(n965) );
  HS65_GS_FA1X4 U959 ( .A0(n875), .B0(n874), .CI(n873), .CO(n878), .S0(n876)
         );
  HS65_GS_IVX2 U960 ( .A(n876), .Z(n958) );
  HS65_GS_FA1X4 U961 ( .A0(n879), .B0(n878), .CI(n877), .CO(n870), .S0(n880)
         );
  HS65_GS_IVX2 U962 ( .A(n880), .Z(n962) );
  HS65_GS_FA1X4 U963 ( .A0(n883), .B0(n882), .CI(n881), .CO(n874), .S0(n884)
         );
  HS65_GS_IVX2 U964 ( .A(n884), .Z(n954) );
  HS65_GS_FA1X4 U965 ( .A0(n887), .B0(n886), .CI(n885), .CO(n882), .S0(n888)
         );
  HS65_GS_IVX2 U966 ( .A(n888), .Z(n950) );
  HS65_GS_FA1X4 U967 ( .A0(n891), .B0(n890), .CI(n889), .CO(n886), .S0(n892)
         );
  HS65_GS_IVX2 U968 ( .A(n892), .Z(n946) );
  HS65_GS_FA1X4 U969 ( .A0(n895), .B0(n894), .CI(n893), .CO(n890), .S0(n896)
         );
  HS65_GS_IVX2 U970 ( .A(n896), .Z(n942) );
  HS65_GS_FA1X4 U971 ( .A0(n899), .B0(n898), .CI(n897), .CO(n894), .S0(n900)
         );
  HS65_GS_IVX2 U972 ( .A(n900), .Z(n938) );
  HS65_GS_FA1X4 U973 ( .A0(n903), .B0(n902), .CI(n901), .CO(n898), .S0(n904)
         );
  HS65_GS_IVX2 U974 ( .A(n904), .Z(n934) );
  HS65_GS_FA1X4 U975 ( .A0(n907), .B0(n906), .CI(n905), .CO(n902), .S0(n908)
         );
  HS65_GS_IVX2 U976 ( .A(n908), .Z(n930) );
  HS65_GS_FA1X4 U977 ( .A0(n911), .B0(n910), .CI(n909), .CO(n906), .S0(n912)
         );
  HS65_GS_IVX2 U978 ( .A(n912), .Z(n926) );
  HS65_GS_FA1X4 U979 ( .A0(n915), .B0(n914), .CI(n913), .CO(n910), .S0(n916)
         );
  HS65_GS_IVX2 U980 ( .A(n916), .Z(n921) );
  HS65_GS_FA1X4 U981 ( .A0(p_b2[1]), .B0(n918), .CI(n917), .CO(n914), .S0(n919) );
  HS65_GS_IVX2 U982 ( .A(n919), .Z(n923) );
  HS65_GS_FA1X4 U983 ( .A0(p_a2[0]), .B0(p_a1[0]), .CI(n920), .CO(n922), .S0(
        n995) );
  HS65_GS_NAND2X2 U984 ( .A(n1335), .B(p_a1[1]), .Z(n1334) );
  HS65_GS_NAND3AX3 U985 ( .A(n1334), .B(p_a2[1]), .C(n923), .Z(n925) );
  HS65_GS_FA1X4 U986 ( .A0(p_a2[2]), .B0(p_a1[2]), .CI(n921), .CO(n928), .S0(
        n1339) );
  HS65_GS_FA1X4 U987 ( .A0(p_a2[1]), .B0(n923), .CI(n922), .CO(n924), .S0(
        n1335) );
  HS65_GS_CB4I1X4 U988 ( .A(p_a1[1]), .B(n1335), .C(n924), .D(n925), .Z(n1338)
         );
  HS65_GS_NAND2X2 U989 ( .A(n1339), .B(n1338), .Z(n1337) );
  HS65_GS_NAND2X2 U990 ( .A(n925), .B(n1337), .Z(n927) );
  HS65_GS_NOR2X2 U991 ( .A(n928), .B(n927), .Z(n929) );
  HS65_GS_FA1X4 U992 ( .A0(p_a2[3]), .B0(p_a1[3]), .CI(n926), .CO(n932), .S0(
        n1343) );
  HS65_GSS_XNOR2X3 U993 ( .A(n928), .B(n927), .Z(n1342) );
  HS65_GS_NOR2X2 U994 ( .A(n1343), .B(n1342), .Z(n1341) );
  HS65_GS_NOR2X2 U995 ( .A(n929), .B(n1341), .Z(n931) );
  HS65_GS_NAND2X2 U996 ( .A(n932), .B(n931), .Z(n933) );
  HS65_GS_FA1X4 U997 ( .A0(p_a2[4]), .B0(p_a1[4]), .CI(n930), .CO(n935), .S0(
        n1347) );
  HS65_GSS_XOR2X3 U998 ( .A(n932), .B(n931), .Z(n1346) );
  HS65_GS_NAND2X2 U999 ( .A(n1347), .B(n1346), .Z(n1345) );
  HS65_GS_NAND2X2 U1000 ( .A(n933), .B(n1345), .Z(n936) );
  HS65_GS_NAND2X2 U1001 ( .A(n935), .B(n936), .Z(n937) );
  HS65_GS_FA1X4 U1002 ( .A0(p_a2[5]), .B0(p_a1[5]), .CI(n934), .CO(n939), .S0(
        n1351) );
  HS65_GSS_XOR2X3 U1003 ( .A(n936), .B(n935), .Z(n1350) );
  HS65_GS_NAND2X2 U1004 ( .A(n1351), .B(n1350), .Z(n1349) );
  HS65_GS_NAND2X2 U1005 ( .A(n937), .B(n1349), .Z(n940) );
  HS65_GS_NAND2X2 U1006 ( .A(n939), .B(n940), .Z(n941) );
  HS65_GS_FA1X4 U1007 ( .A0(p_a2[6]), .B0(p_a1[6]), .CI(n938), .CO(n943), .S0(
        n1355) );
  HS65_GSS_XOR2X3 U1008 ( .A(n940), .B(n939), .Z(n1354) );
  HS65_GS_NAND2X2 U1009 ( .A(n1355), .B(n1354), .Z(n1353) );
  HS65_GS_NAND2X2 U1010 ( .A(n941), .B(n1353), .Z(n944) );
  HS65_GS_NAND2X2 U1011 ( .A(n943), .B(n944), .Z(n945) );
  HS65_GS_FA1X4 U1012 ( .A0(p_a2[7]), .B0(p_a1[7]), .CI(n942), .CO(n947), .S0(
        n1359) );
  HS65_GSS_XOR2X3 U1013 ( .A(n944), .B(n943), .Z(n1358) );
  HS65_GS_NAND2X2 U1014 ( .A(n1359), .B(n1358), .Z(n1357) );
  HS65_GS_NAND2X2 U1015 ( .A(n945), .B(n1357), .Z(n948) );
  HS65_GS_NAND2X2 U1016 ( .A(n947), .B(n948), .Z(n949) );
  HS65_GS_FA1X4 U1017 ( .A0(p_a2[8]), .B0(p_a1[8]), .CI(n946), .CO(n951), .S0(
        n1363) );
  HS65_GSS_XOR2X3 U1018 ( .A(n948), .B(n947), .Z(n1362) );
  HS65_GS_NAND2X2 U1019 ( .A(n1363), .B(n1362), .Z(n1361) );
  HS65_GS_NAND2X2 U1020 ( .A(n949), .B(n1361), .Z(n952) );
  HS65_GS_NAND2X2 U1021 ( .A(n951), .B(n952), .Z(n953) );
  HS65_GS_FA1X4 U1022 ( .A0(p_a2[9]), .B0(p_a1[9]), .CI(n950), .CO(n955), .S0(
        n1367) );
  HS65_GSS_XOR2X3 U1023 ( .A(n952), .B(n951), .Z(n1366) );
  HS65_GS_NAND2X2 U1024 ( .A(n1367), .B(n1366), .Z(n1365) );
  HS65_GS_NAND2X2 U1025 ( .A(n953), .B(n1365), .Z(n956) );
  HS65_GS_NAND2X2 U1026 ( .A(n955), .B(n956), .Z(n957) );
  HS65_GS_FA1X4 U1027 ( .A0(p_a2[10]), .B0(p_a1[10]), .CI(n954), .CO(n959), 
        .S0(n1371) );
  HS65_GSS_XOR2X3 U1028 ( .A(n956), .B(n955), .Z(n1370) );
  HS65_GS_NAND2X2 U1029 ( .A(n1371), .B(n1370), .Z(n1369) );
  HS65_GS_NAND2X2 U1030 ( .A(n957), .B(n1369), .Z(n960) );
  HS65_GS_NAND2X2 U1031 ( .A(n959), .B(n960), .Z(n961) );
  HS65_GS_FA1X4 U1032 ( .A0(p_a2[11]), .B0(p_a1[11]), .CI(n958), .CO(n1377), 
        .S0(n1375) );
  HS65_GSS_XOR2X3 U1033 ( .A(n960), .B(n959), .Z(n1374) );
  HS65_GS_NAND2X2 U1034 ( .A(n1375), .B(n1374), .Z(n1373) );
  HS65_GS_NAND2X2 U1035 ( .A(n961), .B(n1373), .Z(n1378) );
  HS65_GS_PAO2X4 U1036 ( .A(n1377), .B(n1380), .P(n1378), .Z(n963) );
  HS65_GS_FA1X4 U1037 ( .A0(p_a2[12]), .B0(p_a1[12]), .CI(n962), .CO(n964), 
        .S0(n1380) );
  HS65_GSS_XOR2X3 U1038 ( .A(n963), .B(n964), .Z(n1388) );
  HS65_GS_AO22X4 U1039 ( .A(n1387), .B(n1388), .C(n964), .D(n963), .Z(n1393)
         );
  HS65_GS_FA1X4 U1040 ( .A0(p_a1[13]), .B0(p_a2[13]), .CI(n965), .CO(n1392), 
        .S0(n1387) );
  HS65_GS_FA1X4 U1041 ( .A0(n968), .B0(n967), .CI(n966), .CO(n974), .S0(n969)
         );
  HS65_GS_IVX2 U1042 ( .A(n969), .Z(n970) );
  HS65_GS_FA1X4 U1043 ( .A0(p_a1[14]), .B0(p_a2[14]), .CI(n970), .CO(n981), 
        .S0(n1391) );
  HS65_GS_FA1X4 U1044 ( .A0(p_a1[15]), .B0(p_a2[15]), .CI(n971), .CO(n986), 
        .S0(n972) );
  HS65_GS_IVX2 U1045 ( .A(n972), .Z(n980) );
  HS65_GS_FA1X4 U1046 ( .A0(n975), .B0(n974), .CI(n973), .CO(n979), .S0(n971)
         );
  HS65_GS_OAI32X2 U1047 ( .A(p_b0[15]), .B(p_b2[15]), .C(p_b1[15]), .D(n977), 
        .E(n976), .Z(n978) );
  HS65_GSS_XNOR2X3 U1048 ( .A(n979), .B(n978), .Z(n983) );
  HS65_GSS_XNOR2X3 U1049 ( .A(n984), .B(n983), .Z(n985) );
  HS65_GS_NAND2X2 U1050 ( .A(n986), .B(n985), .Z(n988) );
  HS65_GS_FA1X4 U1051 ( .A0(n982), .B0(n981), .CI(n980), .CO(n984), .S0(n993)
         );
  HS65_GS_NAND2X2 U1052 ( .A(n984), .B(n983), .Z(n987) );
  HS65_GS_IVX2 U1053 ( .A(valid_T3), .Z(n1884) );
  HS65_GS_NOR2X2 U1054 ( .A(n986), .B(n985), .Z(n990) );
  HS65_GS_NOR3AX2 U1055 ( .A(n987), .B(n1884), .C(n990), .Z(n1882) );
  HS65_GS_IVX2 U1056 ( .A(n1882), .Z(n991) );
  HS65_GS_AOI12X2 U1057 ( .A(n988), .B(n993), .C(n991), .Z(n1394) );
  HS65_GS_IVX2 U1058 ( .A(n1394), .Z(n1384) );
  HS65_GS_IVX2 U1059 ( .A(n988), .Z(n989) );
  HS65_GS_OAI21X2 U1060 ( .A(n990), .B(n989), .C(valid_T3), .Z(n992) );
  HS65_GS_OAI12X3 U1061 ( .A(n993), .B(n992), .C(n991), .Z(n1385) );
  HS65_GS_IVX2 U1062 ( .A(n1385), .Z(n1397) );
  HS65_GS_NAND2X2 U1063 ( .A(data_out[0]), .B(n1884), .Z(n994) );
  HS65_GS_CBI4I1X3 U1064 ( .A(n995), .B(n1384), .C(n1397), .D(n994), .Z(n1986)
         );
  HS65_GS_MUX21I1X3 U1065 ( .D0(n1492), .D1(data_in[15]), .S0(valid_in), .Z(
        n1893) );
  HS65_GS_MUXI21X2 U1066 ( .D0(n998), .D1(n997), .S0(n996), .Z(n1020) );
  HS65_GS_FA1X4 U1067 ( .A0(n1001), .B0(n1000), .CI(n999), .CO(n1008), .S0(
        n1002) );
  HS65_GS_IVX2 U1068 ( .A(n1002), .Z(n1016) );
  HS65_GS_FA1X4 U1069 ( .A0(n1005), .B0(n1004), .CI(n1003), .CO(n1010), .S0(
        n1015) );
  HS65_GS_FA1X4 U1070 ( .A0(n1008), .B0(n1007), .CI(n1006), .CO(n218), .S0(
        n1014) );
  HS65_GS_FA1X4 U1071 ( .A0(n1011), .B0(n1010), .CI(n1009), .CO(n1001), .S0(
        n1013) );
  HS65_GS_NAND3X2 U1072 ( .A(n1015), .B(n1014), .C(n1013), .Z(n1012) );
  HS65_GS_OAI12X3 U1073 ( .A(n1016), .B(n1012), .C(\mul_b1/result_sat[15] ), 
        .Z(n1878) );
  HS65_GS_OAI21X2 U1074 ( .A(n1019), .B(n1020), .C(n1878), .Z(n1018) );
  HS65_GS_NOR3X1 U1075 ( .A(n1015), .B(n1014), .C(n1013), .Z(n1017) );
  HS65_GS_AOI12X3 U1076 ( .A(n1017), .B(n1016), .C(\mul_b1/result_sat[15] ), 
        .Z(n1483) );
  HS65_GS_IVX2 U1077 ( .A(n1483), .Z(n1880) );
  HS65_GS_CBI4I1X3 U1078 ( .A(n1020), .B(n1019), .C(n1018), .D(n1880), .Z(
        \mul_b1/result_sat[13] ) );
  HS65_GS_IVX2 U1079 ( .A(n1492), .Z(n1891) );
  HS65_GS_IVX2 U1080 ( .A(n1021), .Z(n1024) );
  HS65_GS_IVX2 U1081 ( .A(n1022), .Z(n1023) );
  HS65_GS_AOI22X1 U1082 ( .A(n1025), .B(n1024), .C(n1026), .D(n1023), .Z(n1040) );
  HS65_GS_AOI12X2 U1083 ( .A(n1028), .B(n1027), .C(n1026), .Z(n1038) );
  HS65_GS_FA1X4 U1084 ( .A0(n1031), .B0(n1030), .CI(n1029), .CO(n1032), .S0(
        n1037) );
  HS65_GS_FA1X4 U1085 ( .A0(n1034), .B0(n1033), .CI(n1032), .CO(n509), .S0(
        n1036) );
  HS65_GS_NAND3X2 U1086 ( .A(n1038), .B(n1037), .C(n1036), .Z(n1035) );
  HS65_GS_OAI21X2 U1087 ( .A(n1040), .B(n1035), .C(\mul_b0/result_sat[15] ), 
        .Z(n1554) );
  HS65_GS_OAI21X2 U1088 ( .A(n1042), .B(n1043), .C(n1554), .Z(n1041) );
  HS65_GS_NOR3X1 U1089 ( .A(n1038), .B(n1037), .C(n1036), .Z(n1039) );
  HS65_GS_AOI12X2 U1090 ( .A(n1040), .B(n1039), .C(\mul_b0/result_sat[15] ), 
        .Z(n1557) );
  HS65_GS_IVX2 U1091 ( .A(n1557), .Z(n1072) );
  HS65_GS_CBI4I1X3 U1092 ( .A(n1043), .B(n1042), .C(n1041), .D(n1072), .Z(
        \mul_b0/result_sat[13] ) );
  HS65_GS_OAI21X2 U1093 ( .A(n1045), .B(n1046), .C(n1554), .Z(n1044) );
  HS65_GS_CBI4I1X3 U1094 ( .A(n1046), .B(n1045), .C(n1044), .D(n1072), .Z(
        \mul_b0/result_sat[12] ) );
  HS65_GSS_XOR2X3 U1095 ( .A(n1048), .B(n1047), .Z(n1051) );
  HS65_GS_OAI21X2 U1096 ( .A(n1050), .B(n1051), .C(n1554), .Z(n1049) );
  HS65_GS_CBI4I1X3 U1097 ( .A(n1051), .B(n1050), .C(n1049), .D(n1072), .Z(
        \mul_b0/result_sat[11] ) );
  HS65_GS_IVX2 U1098 ( .A(n1554), .Z(n1556) );
  HS65_GS_AO112X4 U1099 ( .A(n1054), .B(n1053), .C(n1556), .D(n1052), .Z(n1055) );
  HS65_GS_NAND2X2 U1100 ( .A(n1072), .B(n1055), .Z(\mul_b0/result_sat[4] ) );
  HS65_GS_AO112X4 U1101 ( .A(n1058), .B(n1057), .C(n1556), .D(n1056), .Z(n1059) );
  HS65_GS_NAND2X2 U1102 ( .A(n1072), .B(n1059), .Z(\mul_b0/result_sat[3] ) );
  HS65_GS_AO112X4 U1103 ( .A(n1062), .B(n1061), .C(n1556), .D(n1060), .Z(n1063) );
  HS65_GS_NAND2X2 U1104 ( .A(n1072), .B(n1063), .Z(\mul_b0/result_sat[2] ) );
  HS65_GS_AO112X4 U1105 ( .A(n1066), .B(n1065), .C(n1556), .D(n1064), .Z(n1067) );
  HS65_GS_NAND2X2 U1106 ( .A(n1072), .B(n1067), .Z(\mul_b0/result_sat[1] ) );
  HS65_GS_AO112X4 U1107 ( .A(n1070), .B(n1069), .C(n1556), .D(n1068), .Z(n1071) );
  HS65_GS_NAND2X2 U1108 ( .A(n1072), .B(n1071), .Z(\mul_b0/result_sat[0] ) );
  HS65_GS_FA1X4 U1109 ( .A0(n1075), .B0(n1074), .CI(n1073), .CO(n1084), .S0(
        n1076) );
  HS65_GS_IVX2 U1110 ( .A(n1076), .Z(n1091) );
  HS65_GS_FA1X4 U1111 ( .A0(n1079), .B0(n1078), .CI(n1077), .CO(n1082), .S0(
        n1089) );
  HS65_GS_FA1X4 U1112 ( .A0(n1082), .B0(n1081), .CI(n1080), .CO(n740), .S0(
        n1088) );
  HS65_GS_FA1X4 U1113 ( .A0(n1085), .B0(n1084), .CI(n1083), .CO(n1078), .S0(
        n1087) );
  HS65_GS_NAND3X2 U1114 ( .A(n1089), .B(n1088), .C(n1087), .Z(n1086) );
  HS65_GS_OAI12X3 U1115 ( .A(n1091), .B(n1086), .C(\mul_a1/result_sat[15] ), 
        .Z(n1579) );
  HS65_GS_OAI21X2 U1116 ( .A(n1094), .B(n1093), .C(n1579), .Z(n1092) );
  HS65_GS_NOR3X1 U1117 ( .A(n1089), .B(n1088), .C(n1087), .Z(n1090) );
  HS65_GS_AOI12X2 U1118 ( .A(n1091), .B(n1090), .C(\mul_a1/result_sat[15] ), 
        .Z(n1581) );
  HS65_GS_IVX2 U1119 ( .A(n1581), .Z(n1868) );
  HS65_GS_CBI4I1X3 U1120 ( .A(n1094), .B(n1093), .C(n1092), .D(n1868), .Z(
        \mul_a1/result_sat[0] ) );
  HS65_GS_OAI21X2 U1121 ( .A(n1096), .B(n1097), .C(n1579), .Z(n1095) );
  HS65_GS_CBI4I1X3 U1122 ( .A(n1097), .B(n1096), .C(n1095), .D(n1868), .Z(
        \mul_a1/result_sat[3] ) );
  HS65_GSS_XNOR2X3 U1123 ( .A(n1099), .B(n1098), .Z(n1102) );
  HS65_GS_OAI21X2 U1124 ( .A(n1101), .B(n1102), .C(n1579), .Z(n1100) );
  HS65_GS_CBI4I1X3 U1125 ( .A(n1102), .B(n1101), .C(n1100), .D(n1868), .Z(
        \mul_a1/result_sat[4] ) );
  HS65_GSS_XNOR2X3 U1126 ( .A(n1104), .B(n1103), .Z(n1107) );
  HS65_GS_OAI21X2 U1127 ( .A(n1106), .B(n1107), .C(n1579), .Z(n1105) );
  HS65_GS_CBI4I1X3 U1128 ( .A(n1107), .B(n1106), .C(n1105), .D(n1868), .Z(
        \mul_a1/result_sat[5] ) );
  HS65_GSS_XNOR2X3 U1129 ( .A(n1109), .B(n1108), .Z(n1112) );
  HS65_GS_OAI21X2 U1130 ( .A(n1111), .B(n1112), .C(n1579), .Z(n1110) );
  HS65_GS_CBI4I1X3 U1131 ( .A(n1112), .B(n1111), .C(n1110), .D(n1868), .Z(
        \mul_a1/result_sat[8] ) );
  HS65_GSS_XNOR2X3 U1132 ( .A(n1114), .B(n1113), .Z(n1116) );
  HS65_GS_AOI12X2 U1133 ( .A(n1117), .B(n1116), .C(n1581), .Z(n1115) );
  HS65_GS_IVX2 U1134 ( .A(n1579), .Z(n1867) );
  HS65_GS_CBI4I6X2 U1135 ( .A(n1117), .B(n1116), .C(n1115), .D(n1867), .Z(
        \mul_a1/result_sat[11] ) );
  HS65_GSS_XOR2X3 U1136 ( .A(n1119), .B(n1118), .Z(n1141) );
  HS65_GS_FA1X4 U1137 ( .A0(n1122), .B0(n1121), .CI(n1120), .CO(n1128), .S0(
        n1123) );
  HS65_GS_IVX2 U1138 ( .A(n1123), .Z(n1138) );
  HS65_GS_FA1X4 U1139 ( .A0(n1126), .B0(n1125), .CI(n1124), .CO(n421), .S0(
        n1136) );
  HS65_GS_FA1X4 U1140 ( .A0(n1129), .B0(n1128), .CI(n1127), .CO(n1131), .S0(
        n1135) );
  HS65_GS_FA1X4 U1141 ( .A0(n1132), .B0(n1131), .CI(n1130), .CO(n1125), .S0(
        n1134) );
  HS65_GS_NAND3X2 U1142 ( .A(n1136), .B(n1135), .C(n1134), .Z(n1133) );
  HS65_GS_OAI12X3 U1143 ( .A(n1138), .B(n1133), .C(\mul_a2/result_sat[15] ), 
        .Z(n1697) );
  HS65_GS_OAI21X2 U1144 ( .A(n1141), .B(n1142), .C(n1697), .Z(n1140) );
  HS65_GS_NOR3X1 U1145 ( .A(n1136), .B(n1135), .C(n1134), .Z(n1137) );
  HS65_GS_AOI12X3 U1146 ( .A(n1138), .B(n1137), .C(\mul_a2/result_sat[15] ), 
        .Z(n1699) );
  HS65_GS_IVX2 U1147 ( .A(n1699), .Z(n1139) );
  HS65_GS_CBI4I1X3 U1148 ( .A(n1142), .B(n1141), .C(n1140), .D(n1139), .Z(
        \mul_a2/result_sat[0] ) );
  HS65_GS_IVX2 U1149 ( .A(n1143), .Z(n1146) );
  HS65_GS_IVX2 U1150 ( .A(n1144), .Z(n1145) );
  HS65_GS_AOI22X1 U1151 ( .A(n1147), .B(n1146), .C(n1148), .D(n1145), .Z(n1162) );
  HS65_GS_AOI12X2 U1152 ( .A(n1150), .B(n1149), .C(n1148), .Z(n1160) );
  HS65_GS_FA1X4 U1153 ( .A0(n1153), .B0(n1152), .CI(n1151), .CO(n1154), .S0(
        n1159) );
  HS65_GS_FA1X4 U1154 ( .A0(n1156), .B0(n1155), .CI(n1154), .CO(n854), .S0(
        n1158) );
  HS65_GS_NOR3X1 U1155 ( .A(n1160), .B(n1159), .C(n1158), .Z(n1157) );
  HS65_GS_AOI12X2 U1156 ( .A(n1162), .B(n1157), .C(\mul_b2/result_sat[15] ), 
        .Z(n1806) );
  HS65_GS_IVX2 U1157 ( .A(n1806), .Z(n1212) );
  HS65_GS_NAND3X2 U1158 ( .A(n1160), .B(n1159), .C(n1158), .Z(n1161) );
  HS65_GS_OAI21X2 U1159 ( .A(n1162), .B(n1161), .C(\mul_b2/result_sat[15] ), 
        .Z(n1807) );
  HS65_GS_IVX2 U1160 ( .A(n1807), .Z(n1799) );
  HS65_GS_AO112X4 U1161 ( .A(n1165), .B(n1164), .C(n1799), .D(n1163), .Z(n1166) );
  HS65_GS_NAND2X2 U1162 ( .A(n1212), .B(n1166), .Z(\mul_b2/result_sat[0] ) );
  HS65_GS_AOI12X2 U1163 ( .A(n1169), .B(n1168), .C(n1806), .Z(n1167) );
  HS65_GS_CBI4I6X2 U1164 ( .A(n1169), .B(n1168), .C(n1167), .D(n1799), .Z(
        \mul_b2/result_sat[1] ) );
  HS65_GS_AOI12X2 U1165 ( .A(n1172), .B(n1171), .C(n1806), .Z(n1170) );
  HS65_GS_CBI4I6X2 U1166 ( .A(n1172), .B(n1171), .C(n1170), .D(n1799), .Z(
        \mul_b2/result_sat[2] ) );
  HS65_GS_AO112X4 U1167 ( .A(n1175), .B(n1174), .C(n1799), .D(n1173), .Z(n1176) );
  HS65_GS_NAND2X2 U1168 ( .A(n1212), .B(n1176), .Z(\mul_b2/result_sat[3] ) );
  HS65_GS_AOI12X2 U1169 ( .A(n1179), .B(n1178), .C(n1806), .Z(n1177) );
  HS65_GS_CBI4I6X2 U1170 ( .A(n1179), .B(n1178), .C(n1177), .D(n1799), .Z(
        \mul_b2/result_sat[4] ) );
  HS65_GS_AO112X4 U1171 ( .A(n1182), .B(n1181), .C(n1799), .D(n1180), .Z(n1183) );
  HS65_GS_NAND2X2 U1172 ( .A(n1212), .B(n1183), .Z(\mul_b2/result_sat[5] ) );
  HS65_GS_AO112X4 U1173 ( .A(n1186), .B(n1185), .C(n1799), .D(n1184), .Z(n1187) );
  HS65_GS_NAND2X2 U1174 ( .A(n1212), .B(n1187), .Z(\mul_b2/result_sat[6] ) );
  HS65_GS_AO112X4 U1175 ( .A(n1190), .B(n1189), .C(n1799), .D(n1188), .Z(n1191) );
  HS65_GS_NAND2X2 U1176 ( .A(n1212), .B(n1191), .Z(\mul_b2/result_sat[7] ) );
  HS65_GS_AO112X4 U1177 ( .A(n1194), .B(n1193), .C(n1799), .D(n1192), .Z(n1195) );
  HS65_GS_NAND2X2 U1178 ( .A(n1212), .B(n1195), .Z(\mul_b2/result_sat[8] ) );
  HS65_GS_AO112X4 U1179 ( .A(n1198), .B(n1197), .C(n1799), .D(n1196), .Z(n1199) );
  HS65_GS_NAND2X2 U1180 ( .A(n1212), .B(n1199), .Z(\mul_b2/result_sat[9] ) );
  HS65_GS_AO112X4 U1181 ( .A(n1202), .B(n1201), .C(n1799), .D(n1200), .Z(n1203) );
  HS65_GS_NAND2X2 U1182 ( .A(n1212), .B(n1203), .Z(\mul_b2/result_sat[10] ) );
  HS65_GS_AO112X4 U1183 ( .A(n1206), .B(n1205), .C(n1799), .D(n1204), .Z(n1207) );
  HS65_GS_NAND2X2 U1184 ( .A(n1212), .B(n1207), .Z(\mul_b2/result_sat[11] ) );
  HS65_GS_AO112X4 U1185 ( .A(n1210), .B(n1209), .C(n1799), .D(n1208), .Z(n1211) );
  HS65_GS_NAND2X2 U1186 ( .A(n1212), .B(n1211), .Z(\mul_b2/result_sat[12] ) );
  HS65_GS_IVX2 U1187 ( .A(x_reg2[0]), .Z(n1848) );
  HS65_GS_IVX2 U1188 ( .A(x_reg2[2]), .Z(n1847) );
  HS65_GS_NOR2X2 U1189 ( .A(n1848), .B(n1847), .Z(\mul_b2/fa1_c0[2] ) );
  HS65_GS_IVX4 U1190 ( .A(n1409), .Z(n1890) );
  HS65_GS_IVX2 U1191 ( .A(x_z1[14]), .Z(n1494) );
  HS65_GS_IVX2 U1192 ( .A(x_z1[13]), .Z(n1496) );
  HS65_GS_IVX2 U1193 ( .A(x_z1[12]), .Z(n1498) );
  HS65_GS_IVX2 U1194 ( .A(x_z1[11]), .Z(n1500) );
  HS65_GS_IVX2 U1195 ( .A(x_z1[10]), .Z(n1503) );
  HS65_GS_IVX2 U1196 ( .A(x_z1[9]), .Z(n1506) );
  HS65_GS_IVX2 U1197 ( .A(x_z1[8]), .Z(n1509) );
  HS65_GS_IVX2 U1198 ( .A(x_z1[7]), .Z(n1512) );
  HS65_GS_IVX2 U1199 ( .A(x_z1[6]), .Z(n1515) );
  HS65_GS_IVX2 U1200 ( .A(x_z1[5]), .Z(n1502) );
  HS65_GS_IVX2 U1201 ( .A(x_z1[4]), .Z(n1505) );
  HS65_GS_IVX2 U1202 ( .A(x_z1[3]), .Z(n1508) );
  HS65_GS_IVX2 U1203 ( .A(x_z1[2]), .Z(n1511) );
  HS65_GS_IVX2 U1204 ( .A(x_z1[1]), .Z(n1514) );
  HS65_GS_IVX2 U1205 ( .A(x_z1[0]), .Z(n1513) );
  HS65_GS_NOR2X2 U1206 ( .A(n1891), .B(n1214), .Z(n1213) );
  HS65_GSS_XNOR2X3 U1207 ( .A(n1213), .B(n1492), .Z(\mul_b0/fa1_s0[31] ) );
  HS65_GSS_XNOR2X3 U1208 ( .A(x_z1[15]), .B(n1214), .Z(n1516) );
  HS65_GSS_XNOR2X3 U1209 ( .A(n1516), .B(n1492), .Z(\mul_b0/fa1_s0[20] ) );
  HS65_GS_NOR2X2 U1210 ( .A(y_z1[15]), .B(n1612), .Z(n1215) );
  HS65_GSS_XNOR2X3 U1211 ( .A(n1215), .B(n1815), .Z(\mul_a1/fa1_s0[27] ) );
  HS65_GS_NOR2X2 U1212 ( .A(y_z2[15]), .B(n1412), .Z(n1216) );
  HS65_GSS_XNOR2X3 U1213 ( .A(n1216), .B(n1398), .Z(\mul_a2/fa1_s2[31] ) );
  HS65_GS_IVX2 U1214 ( .A(x_z2[14]), .Z(n1773) );
  HS65_GS_IVX2 U1215 ( .A(x_z2[13]), .Z(n1771) );
  HS65_GS_IVX2 U1216 ( .A(x_z2[12]), .Z(n1769) );
  HS65_GS_IVX2 U1217 ( .A(x_z2[11]), .Z(n1767) );
  HS65_GS_IVX2 U1218 ( .A(x_z2[10]), .Z(n1765) );
  HS65_GS_IVX2 U1219 ( .A(x_z2[9]), .Z(n1764) );
  HS65_GS_IVX2 U1220 ( .A(x_z2[8]), .Z(n1760) );
  HS65_GS_IVX2 U1221 ( .A(x_z2[7]), .Z(n1758) );
  HS65_GS_IVX2 U1222 ( .A(x_z2[6]), .Z(n1756) );
  HS65_GS_IVX2 U1223 ( .A(x_z2[5]), .Z(n1763) );
  HS65_GS_IVX2 U1224 ( .A(x_z2[4]), .Z(n1738) );
  HS65_GS_IVX2 U1225 ( .A(x_z2[3]), .Z(n1742) );
  HS65_GS_IVX2 U1226 ( .A(x_z2[2]), .Z(n1747) );
  HS65_GS_IVX2 U1227 ( .A(x_z2[1]), .Z(n1750) );
  HS65_GS_IVX2 U1228 ( .A(x_z2[0]), .Z(n1749) );
  HS65_GS_NOR2X2 U1229 ( .A(x_z2[15]), .B(n1780), .Z(n1217) );
  HS65_GSS_XNOR2X3 U1230 ( .A(n1217), .B(n1810), .Z(\mul_b1/fa1_s0[27] ) );
  HS65_GS_BFX4 U1231 ( .A(valid_in), .Z(n1411) );
  HS65_GS_MUXI21X2 U1232 ( .D0(n1314), .D1(n1842), .S0(n1411), .Z(n1988) );
  HS65_GS_HA1X4 U1233 ( .A0(n1844), .B0(n1314), .CO(n1268), .S0(n1700) );
  HS65_GS_AND2X4 U1234 ( .A(n1700), .B(\mul_a2/fa1_s0[0] ), .Z(
        \mul_a2/fa1_c2[14] ) );
  HS65_GSS_XNOR2X3 U1235 ( .A(n2), .B(n1398), .Z(n1223) );
  HS65_GS_HA1X4 U1236 ( .A0(n1398), .B0(n1218), .CO(n1220), .S0(n1888) );
  HS65_GS_OR2X4 U1237 ( .A(y_z2[15]), .B(n1220), .Z(n1219) );
  HS65_GSS_XNOR2X3 U1238 ( .A(n1223), .B(n1219), .Z(\mul_a2/fa1_s0[27] ) );
  HS65_GSS_XOR2X3 U1239 ( .A(y_z2[15]), .B(n1220), .Z(n1221) );
  HS65_GSS_XNOR2X3 U1240 ( .A(n1223), .B(n1221), .Z(\mul_a2/fa1_s0[20] ) );
  HS65_GS_IVX2 U1241 ( .A(n1888), .Z(n1222) );
  HS65_GSS_XNOR2X3 U1242 ( .A(n1223), .B(n1222), .Z(\mul_a2/fa1_s0[19] ) );
  HS65_GSS_XNOR2X3 U1243 ( .A(y_z2[15]), .B(n1224), .Z(n1253) );
  HS65_GS_HA1X4 U1244 ( .A0(n1726), .B0(n1225), .CO(n1218), .S0(n1252) );
  HS65_GSS_XOR3X2 U1245 ( .A(y_z2[15]), .B(n1253), .C(n1252), .Z(
        \mul_a2/fa1_s0[18] ) );
  HS65_GS_HA1X4 U1246 ( .A0(n1724), .B0(n1226), .CO(n1225), .S0(n1255) );
  HS65_GS_HA1X4 U1247 ( .A0(n1398), .B0(n1227), .CO(n1224), .S0(n1254) );
  HS65_GSS_XOR3X2 U1248 ( .A(y_z2[15]), .B(n1255), .C(n1254), .Z(
        \mul_a2/fa1_s0[17] ) );
  HS65_GS_HA1X4 U1249 ( .A0(n1722), .B0(n1228), .CO(n1226), .S0(n1257) );
  HS65_GS_HA1X4 U1250 ( .A0(n1726), .B0(n1229), .CO(n1227), .S0(n1256) );
  HS65_GSS_XOR3X2 U1251 ( .A(y_z2[15]), .B(n1257), .C(n1256), .Z(
        \mul_a2/fa1_s0[16] ) );
  HS65_GS_HA1X4 U1252 ( .A0(n1720), .B0(n1230), .CO(n1228), .S0(n1259) );
  HS65_GS_HA1X4 U1253 ( .A0(n1724), .B0(n1231), .CO(n1229), .S0(n1258) );
  HS65_GSS_XOR3X2 U1254 ( .A(y_z2[15]), .B(n1259), .C(n1258), .Z(
        \mul_a2/fa1_s0[15] ) );
  HS65_GS_HA1X4 U1255 ( .A0(n1722), .B0(n1232), .CO(n1231), .S0(n1261) );
  HS65_GS_HA1X4 U1256 ( .A0(n1718), .B0(n1233), .CO(n1230), .S0(n1260) );
  HS65_GSS_XOR3X2 U1257 ( .A(y_z2[14]), .B(n1261), .C(n1260), .Z(
        \mul_a2/fa1_s0[14] ) );
  HS65_GS_HA1X4 U1258 ( .A0(n1716), .B0(n1234), .CO(n1233), .S0(n1263) );
  HS65_GS_HA1X4 U1259 ( .A0(n1720), .B0(n1235), .CO(n1232), .S0(n1262) );
  HS65_GSS_XOR3X2 U1260 ( .A(y_z2[13]), .B(n1263), .C(n1262), .Z(
        \mul_a2/fa1_s0[13] ) );
  HS65_GS_HA1X4 U1261 ( .A0(n1718), .B0(n1236), .CO(n1235), .S0(n1265) );
  HS65_GS_HA1X4 U1262 ( .A0(n1714), .B0(n1237), .CO(n1234), .S0(n1264) );
  HS65_GSS_XOR3X2 U1263 ( .A(y_z2[12]), .B(n1265), .C(n1264), .Z(
        \mul_a2/fa1_s0[12] ) );
  HS65_GS_HA1X4 U1264 ( .A0(n1716), .B0(n1238), .CO(n1236), .S0(n1267) );
  HS65_GS_HA1X4 U1265 ( .A0(n1712), .B0(n1239), .CO(n1237), .S0(n1266) );
  HS65_GSS_XOR3X2 U1266 ( .A(y_z2[11]), .B(n1267), .C(n1266), .Z(
        \mul_a2/fa1_s0[11] ) );
  HS65_GS_HA1X4 U1267 ( .A0(n1714), .B0(n1240), .CO(n1238), .S0(n1270) );
  HS65_GS_HA1X4 U1268 ( .A0(n1710), .B0(n1241), .CO(n1239), .S0(n1269) );
  HS65_GSS_XOR3X2 U1269 ( .A(y_z2[10]), .B(n1270), .C(n1269), .Z(
        \mul_a2/fa1_s0[10] ) );
  HS65_GS_HA1X4 U1270 ( .A0(n1712), .B0(n1242), .CO(n1240), .S0(n1272) );
  HS65_GS_HA1X4 U1271 ( .A0(n1708), .B0(n1243), .CO(n1241), .S0(n1271) );
  HS65_GSS_XOR3X2 U1272 ( .A(y_z2[9]), .B(n1272), .C(n1271), .Z(
        \mul_a2/fa1_s0[9] ) );
  HS65_GS_HA1X4 U1273 ( .A0(n1710), .B0(n1244), .CO(n1242), .S0(n1274) );
  HS65_GS_HA1X4 U1274 ( .A0(n1706), .B0(n1245), .CO(n1243), .S0(n1273) );
  HS65_GSS_XOR3X2 U1275 ( .A(y_z2[8]), .B(n1274), .C(n1273), .Z(
        \mul_a2/fa1_s0[8] ) );
  HS65_GS_HA1X4 U1276 ( .A0(n1708), .B0(n1246), .CO(n1244), .S0(n1276) );
  HS65_GS_HA1X4 U1277 ( .A0(n1704), .B0(n1247), .CO(n1245), .S0(n1275) );
  HS65_GSS_XOR3X2 U1278 ( .A(y_z2[7]), .B(n1276), .C(n1275), .Z(
        \mul_a2/fa1_s0[7] ) );
  HS65_GS_HA1X4 U1279 ( .A0(n1706), .B0(n1248), .CO(n1246), .S0(n1278) );
  HS65_GS_HA1X4 U1280 ( .A0(n1702), .B0(n1249), .CO(n1247), .S0(n1277) );
  HS65_GSS_XOR3X2 U1281 ( .A(y_z2[6]), .B(n1278), .C(n1277), .Z(
        \mul_a2/fa1_s0[6] ) );
  HS65_GS_HA1X4 U1282 ( .A0(n1704), .B0(n1250), .CO(n1248), .S0(n1280) );
  HS65_GS_HA1X4 U1283 ( .A0(n1844), .B0(n1314), .CO(n1249), .S0(n1279) );
  HS65_GSS_XOR3X2 U1284 ( .A(y_z2[5]), .B(n1280), .C(n1279), .Z(
        \mul_a2/fa1_s0[5] ) );
  HS65_GS_HA1X4 U1285 ( .A0(n1702), .B0(n1251), .CO(n1250), .S0(n1281) );
  HS65_GSS_XOR3X2 U1286 ( .A(y_z2[4]), .B(n1281), .C(\mul_a2/fa1_s0[0] ), .Z(
        \mul_a2/fa1_s0[4] ) );
  HS65_GS_HA1X4 U1287 ( .A0(n1844), .B0(n1314), .CO(n1251), .S0(n1812) );
  HS65_GSS_XOR2X3 U1288 ( .A(n1812), .B(y_z2[3]), .Z(\mul_a2/fa1_s0[3] ) );
  HS65_GS_PAO2X4 U1289 ( .A(n1253), .B(n1252), .P(y_z2[15]), .Z(
        \mul_a2/fa1_c0[18] ) );
  HS65_GS_PAO2X4 U1290 ( .A(n1255), .B(n1254), .P(y_z2[15]), .Z(
        \mul_a2/fa1_c0[17] ) );
  HS65_GS_PAO2X4 U1291 ( .A(n1257), .B(n1256), .P(y_z2[15]), .Z(
        \mul_a2/fa1_c0[16] ) );
  HS65_GS_PAO2X4 U1292 ( .A(n1259), .B(n1258), .P(y_z2[15]), .Z(
        \mul_a2/fa1_c0[15] ) );
  HS65_GS_PAO2X4 U1293 ( .A(n1261), .B(n1260), .P(y_z2[14]), .Z(
        \mul_a2/fa1_c0[14] ) );
  HS65_GS_PAO2X4 U1294 ( .A(n1263), .B(n1262), .P(y_z2[13]), .Z(
        \mul_a2/fa1_c0[13] ) );
  HS65_GS_PAO2X4 U1295 ( .A(n1265), .B(n1264), .P(y_z2[12]), .Z(
        \mul_a2/fa1_c0[12] ) );
  HS65_GS_PAO2X4 U1296 ( .A(n1267), .B(n1266), .P(y_z2[11]), .Z(
        \mul_a2/fa1_c0[11] ) );
  HS65_GS_HA1X4 U1297 ( .A0(n1702), .B0(n1268), .CO(n1424), .S0(n1701) );
  HS65_GS_AND2X4 U1298 ( .A(n1701), .B(\mul_a2/fa1_s0[1] ), .Z(
        \mul_a2/fa1_c2[15] ) );
  HS65_GS_PAO2X4 U1299 ( .A(n1270), .B(n1269), .P(y_z2[10]), .Z(
        \mul_a2/fa1_c0[10] ) );
  HS65_GS_PAO2X4 U1300 ( .A(n1272), .B(n1271), .P(y_z2[9]), .Z(
        \mul_a2/fa1_c0[9] ) );
  HS65_GS_PAO2X4 U1301 ( .A(n1274), .B(n1273), .P(y_z2[8]), .Z(
        \mul_a2/fa1_c0[8] ) );
  HS65_GS_PAO2X4 U1302 ( .A(n1276), .B(n1275), .P(y_z2[7]), .Z(
        \mul_a2/fa1_c0[7] ) );
  HS65_GS_PAO2X4 U1303 ( .A(n1278), .B(n1277), .P(y_z2[6]), .Z(
        \mul_a2/fa1_c0[6] ) );
  HS65_GS_PAO2X4 U1304 ( .A(n1280), .B(n1279), .P(y_z2[5]), .Z(
        \mul_a2/fa1_c0[5] ) );
  HS65_GS_PAO2X4 U1305 ( .A(n1281), .B(\mul_a2/fa1_s0[0] ), .P(y_z2[4]), .Z(
        \mul_a2/fa1_c0[4] ) );
  HS65_GS_NOR2X2 U1306 ( .A(y_z2[15]), .B(n1283), .Z(n1282) );
  HS65_GSS_XOR3X2 U1307 ( .A(y_z2[15]), .B(n1282), .C(n1), .Z(
        \mul_a2/fa1_s1[27] ) );
  HS65_GSS_XNOR2X3 U1308 ( .A(y_z2[15]), .B(n1283), .Z(n1284) );
  HS65_GSS_XOR3X2 U1309 ( .A(n1), .B(n1284), .C(y_z2[14]), .Z(
        \mul_a2/fa1_s1[24] ) );
  HS65_GS_HA1X4 U1310 ( .A0(n1398), .B0(n1285), .CO(n1283), .S0(n1286) );
  HS65_GSS_XOR3X2 U1311 ( .A(n1), .B(y_z2[13]), .C(n1286), .Z(
        \mul_a2/fa1_s1[23] ) );
  HS65_GSS_XNOR2X3 U1312 ( .A(y_z2[15]), .B(n1287), .Z(n1317) );
  HS65_GS_HA1X4 U1313 ( .A0(n1726), .B0(n1288), .CO(n1285), .S0(n1316) );
  HS65_GSS_XOR3X2 U1314 ( .A(n1317), .B(y_z2[12]), .C(n1316), .Z(
        \mul_a2/fa1_s1[22] ) );
  HS65_GS_HA1X4 U1315 ( .A0(n1724), .B0(n1289), .CO(n1288), .S0(n1319) );
  HS65_GS_HA1X4 U1316 ( .A0(n1398), .B0(n1290), .CO(n1287), .S0(n1318) );
  HS65_GSS_XOR3X2 U1317 ( .A(y_z2[11]), .B(n1319), .C(n1318), .Z(
        \mul_a2/fa1_s1[21] ) );
  HS65_GS_HA1X4 U1318 ( .A0(n1726), .B0(n1291), .CO(n1290), .S0(n1321) );
  HS65_GS_HA1X4 U1319 ( .A0(n1722), .B0(n1292), .CO(n1289), .S0(n1320) );
  HS65_GSS_XOR3X2 U1320 ( .A(y_z2[10]), .B(n1321), .C(n1320), .Z(
        \mul_a2/fa1_s1[20] ) );
  HS65_GS_HA1X4 U1321 ( .A0(n1724), .B0(n1293), .CO(n1291), .S0(n1323) );
  HS65_GS_HA1X4 U1322 ( .A0(n1720), .B0(n1294), .CO(n1292), .S0(n1322) );
  HS65_GSS_XOR3X2 U1323 ( .A(y_z2[9]), .B(n1323), .C(n1322), .Z(
        \mul_a2/fa1_s1[19] ) );
  HS65_GS_HA1X4 U1324 ( .A0(n1722), .B0(n1295), .CO(n1293), .S0(n1325) );
  HS65_GS_HA1X4 U1325 ( .A0(n1718), .B0(n1296), .CO(n1294), .S0(n1324) );
  HS65_GSS_XOR3X2 U1326 ( .A(y_z2[8]), .B(n1325), .C(n1324), .Z(
        \mul_a2/fa1_s1[18] ) );
  HS65_GS_HA1X4 U1327 ( .A0(n1720), .B0(n1297), .CO(n1295), .S0(n1327) );
  HS65_GS_HA1X4 U1328 ( .A0(n1716), .B0(n1298), .CO(n1296), .S0(n1326) );
  HS65_GSS_XOR3X2 U1329 ( .A(y_z2[7]), .B(n1327), .C(n1326), .Z(
        \mul_a2/fa1_s1[17] ) );
  HS65_GS_HA1X4 U1330 ( .A0(n1718), .B0(n1299), .CO(n1297), .S0(n1329) );
  HS65_GS_HA1X4 U1331 ( .A0(n1714), .B0(n1300), .CO(n1298), .S0(n1328) );
  HS65_GSS_XOR3X2 U1332 ( .A(y_z2[6]), .B(n1329), .C(n1328), .Z(
        \mul_a2/fa1_s1[16] ) );
  HS65_GS_HA1X4 U1333 ( .A0(n1716), .B0(n1301), .CO(n1299), .S0(n1331) );
  HS65_GS_HA1X4 U1334 ( .A0(n1712), .B0(n1302), .CO(n1300), .S0(n1330) );
  HS65_GSS_XOR3X2 U1335 ( .A(y_z2[5]), .B(n1331), .C(n1330), .Z(
        \mul_a2/fa1_s1[15] ) );
  HS65_GS_HA1X4 U1336 ( .A0(n1714), .B0(n1303), .CO(n1301), .S0(n1333) );
  HS65_GS_HA1X4 U1337 ( .A0(n1710), .B0(n1304), .CO(n1302), .S0(n1332) );
  HS65_GSS_XOR3X2 U1338 ( .A(y_z2[4]), .B(n1333), .C(n1332), .Z(
        \mul_a2/fa1_s1[14] ) );
  HS65_GS_HA1X4 U1339 ( .A0(n1712), .B0(n1305), .CO(n1303), .S0(n1426) );
  HS65_GS_HA1X4 U1340 ( .A0(n1708), .B0(n1306), .CO(n1304), .S0(n1425) );
  HS65_GSS_XOR3X2 U1341 ( .A(y_z2[3]), .B(n1426), .C(n1425), .Z(
        \mul_a2/fa1_s1[13] ) );
  HS65_GS_HA1X4 U1342 ( .A0(n1706), .B0(n1307), .CO(n1306), .S0(n1736) );
  HS65_GS_HA1X4 U1343 ( .A0(n1710), .B0(n1308), .CO(n1305), .S0(n1735) );
  HS65_GSS_XOR3X2 U1344 ( .A(y_z2[2]), .B(n1736), .C(n1735), .Z(
        \mul_a2/fa1_s1[12] ) );
  HS65_GS_HA1X4 U1345 ( .A0(n1708), .B0(n1309), .CO(n1308), .S0(n1734) );
  HS65_GS_HA1X4 U1346 ( .A0(n1704), .B0(n1310), .CO(n1307), .S0(n1733) );
  HS65_GSS_XOR3X2 U1347 ( .A(\mul_a2/fa1_s0[1] ), .B(n1734), .C(n1733), .Z(
        \mul_a2/fa1_s1[11] ) );
  HS65_GS_HA1X4 U1348 ( .A0(n1706), .B0(n1311), .CO(n1309), .S0(n1732) );
  HS65_GS_HA1X4 U1349 ( .A0(n1702), .B0(n1312), .CO(n1310), .S0(n1731) );
  HS65_GSS_XOR3X2 U1350 ( .A(\mul_a2/fa1_s0[0] ), .B(n1732), .C(n1731), .Z(
        \mul_a2/fa1_s1[10] ) );
  HS65_GS_HA1X4 U1351 ( .A0(n1704), .B0(n1313), .CO(n1311), .S0(n1730) );
  HS65_GS_HA1X4 U1352 ( .A0(n1844), .B0(n1314), .CO(n1312), .S0(n1729) );
  HS65_GSS_XOR2X3 U1353 ( .A(n1730), .B(n1729), .Z(\mul_a2/fa1_s1[9] ) );
  HS65_GS_HA1X4 U1354 ( .A0(n1702), .B0(n1315), .CO(n1313), .S0(n1728) );
  HS65_GSS_XOR2X3 U1355 ( .A(n1728), .B(\mul_a2/fa1_s0[0] ), .Z(
        \mul_a2/fa1_s1[8] ) );
  HS65_GS_PAO2X4 U1356 ( .A(n1317), .B(n1316), .P(y_z2[12]), .Z(
        \mul_a2/fa1_c1[22] ) );
  HS65_GS_PAO2X4 U1357 ( .A(n1319), .B(n1318), .P(y_z2[11]), .Z(
        \mul_a2/fa1_c1[21] ) );
  HS65_GS_PAO2X4 U1358 ( .A(n1321), .B(n1320), .P(y_z2[10]), .Z(
        \mul_a2/fa1_c1[20] ) );
  HS65_GS_PAO2X4 U1359 ( .A(n1323), .B(n1322), .P(y_z2[9]), .Z(
        \mul_a2/fa1_c1[19] ) );
  HS65_GS_PAO2X4 U1360 ( .A(n1325), .B(n1324), .P(y_z2[8]), .Z(
        \mul_a2/fa1_c1[18] ) );
  HS65_GS_PAO2X4 U1361 ( .A(n1327), .B(n1326), .P(y_z2[7]), .Z(
        \mul_a2/fa1_c1[17] ) );
  HS65_GS_PAO2X4 U1362 ( .A(n1329), .B(n1328), .P(y_z2[6]), .Z(
        \mul_a2/fa1_c1[16] ) );
  HS65_GS_PAO2X4 U1363 ( .A(n1331), .B(n1330), .P(y_z2[5]), .Z(
        \mul_a2/fa1_c1[15] ) );
  HS65_GS_PAO2X4 U1364 ( .A(n1333), .B(n1332), .P(y_z2[4]), .Z(
        \mul_a2/fa1_c1[14] ) );
  HS65_GS_MUX21X4 U1365 ( .D0(y_z1[0]), .D1(data_out[0]), .S0(n1892), .Z(n1987) );
  HS65_GS_MUXI21X2 U1366 ( .D0(n1844), .D1(n1843), .S0(n1411), .Z(n1985) );
  HS65_GS_MUX21X4 U1367 ( .D0(y_z1[1]), .D1(data_out[1]), .S0(n1892), .Z(n1984) );
  HS65_GS_OAI112X1 U1368 ( .A(n1335), .B(p_a1[1]), .C(n1384), .D(n1334), .Z(
        n1336) );
  HS65_GS_AO22X4 U1369 ( .A(data_out[1]), .B(n1884), .C(n1385), .D(n1336), .Z(
        n1983) );
  HS65_GS_MUXI21X2 U1370 ( .D0(n1702), .D1(n1841), .S0(n1411), .Z(n1982) );
  HS65_GS_MUX21X4 U1371 ( .D0(y_z1[2]), .D1(data_out[2]), .S0(n1892), .Z(n1981) );
  HS65_GS_OAI112X1 U1372 ( .A(n1339), .B(n1338), .C(n1384), .D(n1337), .Z(
        n1340) );
  HS65_GS_AO22X4 U1373 ( .A(data_out[2]), .B(n1884), .C(n1385), .D(n1340), .Z(
        n1980) );
  HS65_GS_BFX4 U1374 ( .A(valid_in), .Z(n1410) );
  HS65_GS_MUXI21X2 U1375 ( .D0(n1704), .D1(n1839), .S0(n1410), .Z(n1979) );
  HS65_GS_MUX21X4 U1376 ( .D0(y_z1[3]), .D1(data_out[3]), .S0(n1892), .Z(n1978) );
  HS65_GS_AOI112X2 U1377 ( .A(n1343), .B(n1342), .C(n1397), .D(n1341), .Z(
        n1344) );
  HS65_GS_AO112X4 U1378 ( .A(data_out[3]), .B(n1884), .C(n1344), .D(n1394), 
        .Z(n1977) );
  HS65_GS_MUXI21X2 U1379 ( .D0(n1706), .D1(n1837), .S0(n1411), .Z(n1976) );
  HS65_GS_MUX21X4 U1380 ( .D0(y_z1[4]), .D1(data_out[4]), .S0(n1892), .Z(n1975) );
  HS65_GS_OAI112X1 U1381 ( .A(n1347), .B(n1346), .C(n1384), .D(n1345), .Z(
        n1348) );
  HS65_GS_AO22X4 U1382 ( .A(data_out[4]), .B(n1884), .C(n1385), .D(n1348), .Z(
        n1974) );
  HS65_GS_MUXI21X2 U1383 ( .D0(n1708), .D1(n1835), .S0(n1411), .Z(n1973) );
  HS65_GS_MUX21X4 U1384 ( .D0(y_z1[5]), .D1(data_out[5]), .S0(valid_in), .Z(
        n1972) );
  HS65_GS_OAI112X1 U1385 ( .A(n1351), .B(n1350), .C(n1384), .D(n1349), .Z(
        n1352) );
  HS65_GS_AO22X4 U1386 ( .A(data_out[5]), .B(n1884), .C(n1385), .D(n1352), .Z(
        n1971) );
  HS65_GS_MUXI21X2 U1387 ( .D0(n1710), .D1(n1833), .S0(n1411), .Z(n1970) );
  HS65_GS_MUX21X4 U1388 ( .D0(y_z1[6]), .D1(data_out[6]), .S0(n1411), .Z(n1969) );
  HS65_GS_OAI112X1 U1389 ( .A(n1355), .B(n1354), .C(n1384), .D(n1353), .Z(
        n1356) );
  HS65_GS_AO22X4 U1390 ( .A(data_out[6]), .B(n1884), .C(n1385), .D(n1356), .Z(
        n1968) );
  HS65_GS_MUXI21X2 U1391 ( .D0(n1712), .D1(n1831), .S0(n1411), .Z(n1967) );
  HS65_GS_MUX21X4 U1392 ( .D0(y_z1[7]), .D1(data_out[7]), .S0(n1892), .Z(n1966) );
  HS65_GS_OAI112X1 U1393 ( .A(n1359), .B(n1358), .C(n1384), .D(n1357), .Z(
        n1360) );
  HS65_GS_AO22X4 U1394 ( .A(data_out[7]), .B(n1884), .C(n1385), .D(n1360), .Z(
        n1965) );
  HS65_GS_MUXI21X2 U1395 ( .D0(n1714), .D1(n1829), .S0(n1411), .Z(n1964) );
  HS65_GS_MUX21X4 U1396 ( .D0(y_z1[8]), .D1(data_out[8]), .S0(valid_in), .Z(
        n1963) );
  HS65_GS_OAI112X1 U1397 ( .A(n1363), .B(n1362), .C(n1384), .D(n1361), .Z(
        n1364) );
  HS65_GS_AO22X4 U1398 ( .A(data_out[8]), .B(n1884), .C(n1385), .D(n1364), .Z(
        n1962) );
  HS65_GS_MUXI21X2 U1399 ( .D0(n1716), .D1(n1827), .S0(n1411), .Z(n1961) );
  HS65_GS_MUX21X4 U1400 ( .D0(y_z1[9]), .D1(data_out[9]), .S0(valid_in), .Z(
        n1960) );
  HS65_GS_OAI112X1 U1401 ( .A(n1367), .B(n1366), .C(n1384), .D(n1365), .Z(
        n1368) );
  HS65_GS_AO22X4 U1402 ( .A(data_out[9]), .B(n1884), .C(n1385), .D(n1368), .Z(
        n1959) );
  HS65_GS_MUXI21X2 U1403 ( .D0(n1718), .D1(n1825), .S0(n1411), .Z(n1958) );
  HS65_GS_MUX21X4 U1404 ( .D0(y_z1[10]), .D1(data_out[10]), .S0(n1892), .Z(
        n1957) );
  HS65_GS_OAI112X1 U1405 ( .A(n1371), .B(n1370), .C(n1384), .D(n1369), .Z(
        n1372) );
  HS65_GS_AO22X4 U1406 ( .A(data_out[10]), .B(n1884), .C(n1385), .D(n1372), 
        .Z(n1956) );
  HS65_GS_MUXI21X2 U1407 ( .D0(n1720), .D1(n1823), .S0(n1411), .Z(n1955) );
  HS65_GS_MUX21X4 U1408 ( .D0(y_z1[11]), .D1(data_out[11]), .S0(valid_in), .Z(
        n1954) );
  HS65_GS_OAI112X1 U1409 ( .A(n1375), .B(n1374), .C(n1384), .D(n1373), .Z(
        n1376) );
  HS65_GS_AO22X4 U1410 ( .A(data_out[11]), .B(n1884), .C(n1385), .D(n1376), 
        .Z(n1953) );
  HS65_GS_MUXI21X2 U1411 ( .D0(n1722), .D1(n1821), .S0(n1411), .Z(n1952) );
  HS65_GS_IVX2 U1412 ( .A(data_out[12]), .Z(n1383) );
  HS65_GS_MUXI21X2 U1413 ( .D0(n1821), .D1(n1383), .S0(n1411), .Z(n1951) );
  HS65_GSS_XOR2X3 U1414 ( .A(n1378), .B(n1377), .Z(n1381) );
  HS65_GS_OAI21X2 U1415 ( .A(n1380), .B(n1381), .C(n1384), .Z(n1379) );
  HS65_GS_CBI4I1X3 U1416 ( .A(n1381), .B(n1380), .C(n1379), .D(n1385), .Z(
        n1382) );
  HS65_GS_OAI21X2 U1417 ( .A(valid_T3), .B(n1383), .C(n1382), .Z(n1950) );
  HS65_GS_MUXI21X2 U1418 ( .D0(n1724), .D1(n1819), .S0(n1410), .Z(n1949) );
  HS65_GS_IVX2 U1419 ( .A(data_out[13]), .Z(n1390) );
  HS65_GS_MUXI21X2 U1420 ( .D0(n1819), .D1(n1390), .S0(n1410), .Z(n1948) );
  HS65_GS_OAI21X2 U1421 ( .A(n1387), .B(n1388), .C(n1384), .Z(n1386) );
  HS65_GS_CBI4I1X3 U1422 ( .A(n1388), .B(n1387), .C(n1386), .D(n1385), .Z(
        n1389) );
  HS65_GS_OAI21X2 U1423 ( .A(valid_T3), .B(n1390), .C(n1389), .Z(n1947) );
  HS65_GS_MUXI21X2 U1424 ( .D0(n1726), .D1(n1817), .S0(n1410), .Z(n1946) );
  HS65_GS_MUX21X4 U1425 ( .D0(y_z1[14]), .D1(data_out[14]), .S0(n1406), .Z(
        n1945) );
  HS65_GS_FA1X4 U1426 ( .A0(n1393), .B0(n1392), .CI(n1391), .CO(n982), .S0(
        n1396) );
  HS65_GS_AOI12X2 U1427 ( .A(data_out[14]), .B(n1884), .C(n1394), .Z(n1395) );
  HS65_GS_OAI21X2 U1428 ( .A(n1397), .B(n1396), .C(n1395), .Z(n1944) );
  HS65_GS_MUXI21X2 U1429 ( .D0(n1398), .D1(n1815), .S0(n1410), .Z(n1943) );
  HS65_GS_IVX2 U1430 ( .A(data_out[15]), .Z(n1883) );
  HS65_GS_MUXI21X2 U1431 ( .D0(n1815), .D1(n1883), .S0(n1410), .Z(n1942) );
  HS65_GS_MUX21X4 U1432 ( .D0(x_reg2[0]), .D1(x_z2[0]), .S0(n1892), .Z(n1940)
         );
  HS65_GS_MUXI21X2 U1433 ( .D0(n1749), .D1(n1513), .S0(valid_in), .Z(n1939) );
  HS65_GS_MUX21X4 U1434 ( .D0(x_reg2[1]), .D1(x_z2[1]), .S0(valid_in), .Z(
        n1938) );
  HS65_GS_MUXI21X2 U1435 ( .D0(n1750), .D1(n1514), .S0(n1411), .Z(n1937) );
  HS65_GS_MUXI21X2 U1436 ( .D0(n1847), .D1(n1747), .S0(valid_in), .Z(n1936) );
  HS65_GS_MUXI21X2 U1437 ( .D0(n1747), .D1(n1511), .S0(n1406), .Z(n1935) );
  HS65_GS_MUXI21X2 U1438 ( .D0(n1845), .D1(n1742), .S0(n1892), .Z(n1934) );
  HS65_GS_MUXI21X2 U1439 ( .D0(n1742), .D1(n1508), .S0(valid_in), .Z(n1933) );
  HS65_GS_IVX2 U1440 ( .A(x_reg2[4]), .Z(n1850) );
  HS65_GS_MUXI21X2 U1441 ( .D0(n1850), .D1(n1738), .S0(valid_in), .Z(n1932) );
  HS65_GS_MUXI21X2 U1442 ( .D0(n1738), .D1(n1505), .S0(n1406), .Z(n1931) );
  HS65_GS_IVX2 U1443 ( .A(x_reg2[5]), .Z(n1851) );
  HS65_GS_MUXI21X2 U1444 ( .D0(n1851), .D1(n1763), .S0(n1892), .Z(n1930) );
  HS65_GS_MUXI21X2 U1445 ( .D0(n1763), .D1(n1502), .S0(valid_in), .Z(n1929) );
  HS65_GS_IVX2 U1446 ( .A(x_reg2[6]), .Z(n1399) );
  HS65_GS_MUXI21X2 U1447 ( .D0(n1399), .D1(n1756), .S0(n1406), .Z(n1928) );
  HS65_GS_MUXI21X2 U1448 ( .D0(n1756), .D1(n1515), .S0(n1406), .Z(n1927) );
  HS65_GS_IVX2 U1449 ( .A(x_reg2[7]), .Z(n1400) );
  HS65_GS_MUXI21X2 U1450 ( .D0(n1400), .D1(n1758), .S0(n1406), .Z(n1926) );
  HS65_GS_MUXI21X2 U1451 ( .D0(n1758), .D1(n1512), .S0(n1406), .Z(n1925) );
  HS65_GS_IVX2 U1452 ( .A(x_reg2[8]), .Z(n1401) );
  HS65_GS_MUXI21X2 U1453 ( .D0(n1401), .D1(n1760), .S0(n1406), .Z(n1924) );
  HS65_GS_MUXI21X2 U1454 ( .D0(n1760), .D1(n1509), .S0(n1406), .Z(n1923) );
  HS65_GS_IVX2 U1455 ( .A(x_reg2[9]), .Z(n1402) );
  HS65_GS_MUXI21X2 U1456 ( .D0(n1402), .D1(n1764), .S0(n1406), .Z(n1922) );
  HS65_GS_MUXI21X2 U1457 ( .D0(n1764), .D1(n1506), .S0(n1406), .Z(n1921) );
  HS65_GS_IVX2 U1458 ( .A(x_reg2[10]), .Z(n1403) );
  HS65_GS_MUXI21X2 U1459 ( .D0(n1403), .D1(n1765), .S0(n1406), .Z(n1920) );
  HS65_GS_MUXI21X2 U1460 ( .D0(n1765), .D1(n1503), .S0(n1406), .Z(n1919) );
  HS65_GS_IVX2 U1461 ( .A(x_reg2[11]), .Z(n1404) );
  HS65_GS_MUXI21X2 U1462 ( .D0(n1404), .D1(n1767), .S0(n1406), .Z(n1918) );
  HS65_GS_MUXI21X2 U1463 ( .D0(n1767), .D1(n1500), .S0(n1406), .Z(n1917) );
  HS65_GS_IVX2 U1464 ( .A(x_reg2[12]), .Z(n1405) );
  HS65_GS_MUXI21X2 U1465 ( .D0(n1405), .D1(n1769), .S0(n1410), .Z(n1916) );
  HS65_GS_MUXI21X2 U1466 ( .D0(n1769), .D1(n1498), .S0(n1406), .Z(n1915) );
  HS65_GS_IVX2 U1467 ( .A(x_reg2[13]), .Z(n1407) );
  HS65_GS_MUXI21X2 U1468 ( .D0(n1407), .D1(n1771), .S0(n1410), .Z(n1914) );
  HS65_GS_MUXI21X2 U1469 ( .D0(n1771), .D1(n1496), .S0(n1410), .Z(n1913) );
  HS65_GS_IVX2 U1470 ( .A(x_reg2[14]), .Z(n1408) );
  HS65_GS_MUXI21X2 U1471 ( .D0(n1408), .D1(n1773), .S0(n1410), .Z(n1912) );
  HS65_GS_MUXI21X2 U1472 ( .D0(n1773), .D1(n1494), .S0(n1410), .Z(n1911) );
  HS65_GS_MUXI21X2 U1473 ( .D0(n1409), .D1(n1810), .S0(n1410), .Z(n1910) );
  HS65_GS_MUXI21X2 U1474 ( .D0(n1810), .D1(n1492), .S0(n1410), .Z(n1909) );
  HS65_GS_MUX21X4 U1475 ( .D0(x_z1[0]), .D1(data_in[0]), .S0(n1892), .Z(n1908)
         );
  HS65_GS_MUX21X4 U1476 ( .D0(x_z1[1]), .D1(data_in[1]), .S0(valid_in), .Z(
        n1907) );
  HS65_GS_MUX21X4 U1477 ( .D0(x_z1[2]), .D1(data_in[2]), .S0(n1892), .Z(n1906)
         );
  HS65_GS_MUX21X4 U1478 ( .D0(x_z1[3]), .D1(data_in[3]), .S0(n1892), .Z(n1905)
         );
  HS65_GS_MUX21X4 U1479 ( .D0(x_z1[4]), .D1(data_in[4]), .S0(n1411), .Z(n1904)
         );
  HS65_GS_MUX21X4 U1480 ( .D0(x_z1[5]), .D1(data_in[5]), .S0(valid_in), .Z(
        n1903) );
  HS65_GS_MUX21X4 U1481 ( .D0(x_z1[6]), .D1(data_in[6]), .S0(n1892), .Z(n1902)
         );
  HS65_GS_MUX21X4 U1482 ( .D0(x_z1[7]), .D1(data_in[7]), .S0(valid_in), .Z(
        n1901) );
  HS65_GS_MUX21X4 U1483 ( .D0(x_z1[8]), .D1(data_in[8]), .S0(valid_in), .Z(
        n1900) );
  HS65_GS_MUX21X4 U1484 ( .D0(x_z1[9]), .D1(data_in[9]), .S0(n1892), .Z(n1899)
         );
  HS65_GS_MUX21X4 U1485 ( .D0(x_z1[10]), .D1(data_in[10]), .S0(n1892), .Z(
        n1898) );
  HS65_GS_MUX21X4 U1486 ( .D0(x_z1[11]), .D1(data_in[11]), .S0(n1411), .Z(
        n1897) );
  HS65_GS_MUX21X4 U1487 ( .D0(x_z1[12]), .D1(data_in[12]), .S0(n1411), .Z(
        n1896) );
  HS65_GS_MUX21X4 U1488 ( .D0(x_z1[13]), .D1(data_in[13]), .S0(n1892), .Z(
        n1895) );
  HS65_GS_MUX21X4 U1489 ( .D0(x_z1[14]), .D1(data_in[14]), .S0(valid_in), .Z(
        n1894) );
  HS65_GSS_XNOR2X3 U1490 ( .A(y_z2[15]), .B(n1412), .Z(n1727) );
  HS65_GS_AND2X4 U1491 ( .A(y_z2[14]), .B(n1727), .Z(\mul_a2/fa1_c2[28] ) );
  HS65_GS_HA1X4 U1492 ( .A0(n1726), .B0(n1413), .CO(n1412), .S0(n1725) );
  HS65_GS_AND2X4 U1493 ( .A(n1725), .B(y_z2[13]), .Z(\mul_a2/fa1_c2[27] ) );
  HS65_GS_HA1X4 U1494 ( .A0(n1724), .B0(n1414), .CO(n1413), .S0(n1723) );
  HS65_GS_AND2X4 U1495 ( .A(y_z2[12]), .B(n1723), .Z(\mul_a2/fa1_c2[26] ) );
  HS65_GS_HA1X4 U1496 ( .A0(n1722), .B0(n1415), .CO(n1414), .S0(n1721) );
  HS65_GS_AND2X4 U1497 ( .A(n1721), .B(y_z2[11]), .Z(\mul_a2/fa1_c2[25] ) );
  HS65_GS_HA1X4 U1498 ( .A0(n1720), .B0(n1416), .CO(n1415), .S0(n1719) );
  HS65_GS_AND2X4 U1499 ( .A(n1719), .B(y_z2[10]), .Z(\mul_a2/fa1_c2[24] ) );
  HS65_GS_HA1X4 U1500 ( .A0(n1718), .B0(n1417), .CO(n1416), .S0(n1717) );
  HS65_GS_AND2X4 U1501 ( .A(n1717), .B(y_z2[9]), .Z(\mul_a2/fa1_c2[23] ) );
  HS65_GS_HA1X4 U1502 ( .A0(n1716), .B0(n1418), .CO(n1417), .S0(n1715) );
  HS65_GS_AND2X4 U1503 ( .A(n1715), .B(y_z2[8]), .Z(\mul_a2/fa1_c2[22] ) );
  HS65_GS_HA1X4 U1504 ( .A0(n1714), .B0(n1419), .CO(n1418), .S0(n1713) );
  HS65_GS_AND2X4 U1505 ( .A(n1713), .B(y_z2[7]), .Z(\mul_a2/fa1_c2[21] ) );
  HS65_GS_HA1X4 U1506 ( .A0(n1712), .B0(n1420), .CO(n1419), .S0(n1711) );
  HS65_GS_AND2X4 U1507 ( .A(n1711), .B(y_z2[6]), .Z(\mul_a2/fa1_c2[20] ) );
  HS65_GS_HA1X4 U1508 ( .A0(n1710), .B0(n1421), .CO(n1420), .S0(n1709) );
  HS65_GS_AND2X4 U1509 ( .A(n1709), .B(y_z2[5]), .Z(\mul_a2/fa1_c2[19] ) );
  HS65_GS_HA1X4 U1510 ( .A0(n1708), .B0(n1422), .CO(n1421), .S0(n1707) );
  HS65_GS_AND2X4 U1511 ( .A(n1707), .B(y_z2[4]), .Z(\mul_a2/fa1_c2[18] ) );
  HS65_GS_HA1X4 U1512 ( .A0(n1706), .B0(n1423), .CO(n1422), .S0(n1705) );
  HS65_GS_AND2X4 U1513 ( .A(n1705), .B(y_z2[3]), .Z(\mul_a2/fa1_c2[17] ) );
  HS65_GS_HA1X4 U1514 ( .A0(n1704), .B0(n1424), .CO(n1423), .S0(n1703) );
  HS65_GS_AND2X4 U1515 ( .A(n1703), .B(y_z2[2]), .Z(\mul_a2/fa1_c2[16] ) );
  HS65_GS_PAO2X4 U1516 ( .A(n1426), .B(n1425), .P(y_z2[3]), .Z(
        \mul_a2/fa1_c1[13] ) );
  HS65_GSS_XNOR2X3 U1517 ( .A(x_z2[15]), .B(n1809), .Z(n1796) );
  HS65_GSS_XNOR2X3 U1518 ( .A(n1796), .B(n1773), .Z(\mul_b1/fa1_s2[28] ) );
  HS65_GS_HA1X4 U1519 ( .A0(n1773), .B0(n1427), .CO(n1809), .S0(n1795) );
  HS65_GSS_XNOR2X3 U1520 ( .A(n1795), .B(n1771), .Z(\mul_b1/fa1_s2[27] ) );
  HS65_GS_HA1X4 U1521 ( .A0(n1771), .B0(n1428), .CO(n1427), .S0(n1794) );
  HS65_GSS_XNOR2X3 U1522 ( .A(n1794), .B(n1769), .Z(\mul_b1/fa1_s2[26] ) );
  HS65_GS_HA1X4 U1523 ( .A0(n1769), .B0(n1429), .CO(n1428), .S0(n1793) );
  HS65_GSS_XNOR2X3 U1524 ( .A(n1793), .B(n1767), .Z(\mul_b1/fa1_s2[25] ) );
  HS65_GS_HA1X4 U1525 ( .A0(n1767), .B0(n1430), .CO(n1429), .S0(n1792) );
  HS65_GSS_XNOR2X3 U1526 ( .A(n1792), .B(n1765), .Z(\mul_b1/fa1_s2[24] ) );
  HS65_GS_HA1X4 U1527 ( .A0(n1765), .B0(n1431), .CO(n1430), .S0(n1791) );
  HS65_GSS_XNOR2X3 U1528 ( .A(n1791), .B(n1764), .Z(\mul_b1/fa1_s2[23] ) );
  HS65_GS_HA1X4 U1529 ( .A0(n1764), .B0(n1432), .CO(n1431), .S0(n1790) );
  HS65_GSS_XNOR2X3 U1530 ( .A(n1790), .B(n1760), .Z(\mul_b1/fa1_s2[22] ) );
  HS65_GS_HA1X4 U1531 ( .A0(n1760), .B0(n1433), .CO(n1432), .S0(n1789) );
  HS65_GSS_XNOR2X3 U1532 ( .A(n1789), .B(n1758), .Z(\mul_b1/fa1_s2[21] ) );
  HS65_GS_HA1X4 U1533 ( .A0(n1758), .B0(n1434), .CO(n1433), .S0(n1788) );
  HS65_GSS_XNOR2X3 U1534 ( .A(n1788), .B(n1756), .Z(\mul_b1/fa1_s2[20] ) );
  HS65_GS_HA1X4 U1535 ( .A0(n1756), .B0(n1435), .CO(n1434), .S0(n1787) );
  HS65_GSS_XNOR2X3 U1536 ( .A(n1787), .B(n1763), .Z(\mul_b1/fa1_s2[19] ) );
  HS65_GS_HA1X4 U1537 ( .A0(n1763), .B0(n1436), .CO(n1435), .S0(n1786) );
  HS65_GSS_XNOR2X3 U1538 ( .A(n1786), .B(n1738), .Z(\mul_b1/fa1_s2[18] ) );
  HS65_GS_HA1X4 U1539 ( .A0(n1738), .B0(n1437), .CO(n1436), .S0(n1785) );
  HS65_GSS_XNOR2X3 U1540 ( .A(n1785), .B(n1742), .Z(\mul_b1/fa1_s2[17] ) );
  HS65_GS_HA1X4 U1541 ( .A0(n1742), .B0(n1438), .CO(n1437), .S0(n1784) );
  HS65_GSS_XNOR2X3 U1542 ( .A(n1784), .B(n1747), .Z(\mul_b1/fa1_s2[16] ) );
  HS65_GS_HA1X4 U1543 ( .A0(n1747), .B0(n1439), .CO(n1438), .S0(n1783) );
  HS65_GSS_XNOR2X3 U1544 ( .A(n1783), .B(n1750), .Z(\mul_b1/fa1_s2[15] ) );
  HS65_GS_HA1X4 U1545 ( .A0(n1750), .B0(n1749), .CO(n1439), .S0(n1782) );
  HS65_GSS_XNOR2X3 U1546 ( .A(n1782), .B(n1749), .Z(\mul_b1/fa1_s2[14] ) );
  HS65_GS_FA1X4 U1547 ( .A0(n1442), .B0(n1441), .CI(n1440), .CO(n997), .S0(
        n1443) );
  HS65_GS_AO12X4 U1548 ( .A(n1443), .B(n1878), .C(n1483), .Z(
        \mul_b1/result_sat[12] ) );
  HS65_GS_FA1X4 U1549 ( .A0(n1446), .B0(n1445), .CI(n1444), .CO(n1440), .S0(
        n1447) );
  HS65_GS_OA12X4 U1550 ( .A(n1483), .B(n1447), .C(n1878), .Z(
        \mul_b1/result_sat[11] ) );
  HS65_GS_FA1X4 U1551 ( .A0(n1450), .B0(n1449), .CI(n1448), .CO(n1445), .S0(
        n1451) );
  HS65_GS_OA12X4 U1552 ( .A(n1483), .B(n1451), .C(n1878), .Z(
        \mul_b1/result_sat[10] ) );
  HS65_GS_FA1X4 U1553 ( .A0(n1454), .B0(n1453), .CI(n1452), .CO(n1449), .S0(
        n1455) );
  HS65_GS_AO12X4 U1554 ( .A(n1455), .B(n1878), .C(n1483), .Z(
        \mul_b1/result_sat[9] ) );
  HS65_GS_FA1X4 U1555 ( .A0(n1458), .B0(n1457), .CI(n1456), .CO(n1454), .S0(
        n1459) );
  HS65_GS_OA12X4 U1556 ( .A(n1483), .B(n1459), .C(n1878), .Z(
        \mul_b1/result_sat[8] ) );
  HS65_GS_FA1X4 U1557 ( .A0(n1462), .B0(n1461), .CI(n1460), .CO(n1457), .S0(
        n1463) );
  HS65_GS_OA12X4 U1558 ( .A(n1483), .B(n1463), .C(n1878), .Z(
        \mul_b1/result_sat[7] ) );
  HS65_GS_FA1X4 U1559 ( .A0(n1466), .B0(n1465), .CI(n1464), .CO(n1461), .S0(
        n1467) );
  HS65_GS_AO12X4 U1560 ( .A(n1467), .B(n1878), .C(n1483), .Z(
        \mul_b1/result_sat[6] ) );
  HS65_GS_FA1X4 U1561 ( .A0(n1470), .B0(n1469), .CI(n1468), .CO(n1466), .S0(
        n1471) );
  HS65_GS_OA12X4 U1562 ( .A(n1483), .B(n1471), .C(n1878), .Z(
        \mul_b1/result_sat[5] ) );
  HS65_GS_FA1X4 U1563 ( .A0(n1474), .B0(n1473), .CI(n1472), .CO(n1469), .S0(
        n1475) );
  HS65_GS_OA12X4 U1564 ( .A(n1483), .B(n1475), .C(n1878), .Z(
        \mul_b1/result_sat[4] ) );
  HS65_GS_FA1X4 U1565 ( .A0(n1477), .B0(n1479), .CI(n1476), .CO(n1473), .S0(
        n1478) );
  HS65_GS_AO12X4 U1566 ( .A(n1478), .B(n1878), .C(n1483), .Z(
        \mul_b1/result_sat[3] ) );
  HS65_GS_AOI12X2 U1567 ( .A(n1481), .B(n1480), .C(n1479), .Z(n1482) );
  HS65_GS_OA12X4 U1568 ( .A(n1483), .B(n1482), .C(n1878), .Z(
        \mul_b1/result_sat[2] ) );
  HS65_GS_OAI21X2 U1569 ( .A(n1484), .B(n1870), .C(n1878), .Z(n1485) );
  HS65_GS_OAI21X2 U1570 ( .A(n1486), .B(n1485), .C(n1880), .Z(
        \mul_b1/result_sat[1] ) );
  HS65_GS_HA1X4 U1571 ( .A0(n1494), .B0(n1487), .CO(n1214), .S0(n1517) );
  HS65_GSS_XNOR2X3 U1572 ( .A(n1517), .B(n1492), .Z(\mul_b0/fa1_s0[19] ) );
  HS65_GS_HA1X4 U1573 ( .A0(n1496), .B0(n1488), .CO(n1487), .S0(n1518) );
  HS65_GSS_XNOR2X3 U1574 ( .A(n1518), .B(n1492), .Z(\mul_b0/fa1_s0[18] ) );
  HS65_GS_HA1X4 U1575 ( .A0(n1498), .B0(n1489), .CO(n1488), .S0(n1519) );
  HS65_GSS_XNOR2X3 U1576 ( .A(n1519), .B(n1492), .Z(\mul_b0/fa1_s0[17] ) );
  HS65_GS_HA1X4 U1577 ( .A0(n1500), .B0(n1490), .CO(n1489), .S0(n1520) );
  HS65_GSS_XNOR2X3 U1578 ( .A(n1520), .B(n1492), .Z(\mul_b0/fa1_s0[16] ) );
  HS65_GS_HA1X4 U1579 ( .A0(n1503), .B0(n1491), .CO(n1490), .S0(n1521) );
  HS65_GSS_XNOR2X3 U1580 ( .A(n1521), .B(n1492), .Z(\mul_b0/fa1_s0[15] ) );
  HS65_GS_HA1X4 U1581 ( .A0(n1506), .B0(n1493), .CO(n1491), .S0(n1522) );
  HS65_GSS_XNOR2X3 U1582 ( .A(n1522), .B(n1494), .Z(\mul_b0/fa1_s0[14] ) );
  HS65_GS_HA1X4 U1583 ( .A0(n1509), .B0(n1495), .CO(n1493), .S0(n1523) );
  HS65_GSS_XNOR2X3 U1584 ( .A(n1523), .B(n1496), .Z(\mul_b0/fa1_s0[13] ) );
  HS65_GS_HA1X4 U1585 ( .A0(n1512), .B0(n1497), .CO(n1495), .S0(n1524) );
  HS65_GSS_XNOR2X3 U1586 ( .A(n1524), .B(n1498), .Z(\mul_b0/fa1_s0[12] ) );
  HS65_GS_HA1X4 U1587 ( .A0(n1515), .B0(n1499), .CO(n1497), .S0(n1525) );
  HS65_GSS_XNOR2X3 U1588 ( .A(n1525), .B(n1500), .Z(\mul_b0/fa1_s0[11] ) );
  HS65_GS_HA1X4 U1589 ( .A0(n1502), .B0(n1501), .CO(n1499), .S0(n1526) );
  HS65_GSS_XNOR2X3 U1590 ( .A(n1526), .B(n1503), .Z(\mul_b0/fa1_s0[10] ) );
  HS65_GS_HA1X4 U1591 ( .A0(n1505), .B0(n1504), .CO(n1501), .S0(n1527) );
  HS65_GSS_XNOR2X3 U1592 ( .A(n1527), .B(n1506), .Z(\mul_b0/fa1_s0[9] ) );
  HS65_GS_HA1X4 U1593 ( .A0(n1508), .B0(n1507), .CO(n1504), .S0(n1528) );
  HS65_GSS_XNOR2X3 U1594 ( .A(n1528), .B(n1509), .Z(\mul_b0/fa1_s0[8] ) );
  HS65_GS_HA1X4 U1595 ( .A0(n1511), .B0(n1510), .CO(n1507), .S0(n1529) );
  HS65_GSS_XNOR2X3 U1596 ( .A(n1529), .B(n1512), .Z(\mul_b0/fa1_s0[7] ) );
  HS65_GS_HA1X4 U1597 ( .A0(n1514), .B0(n1513), .CO(n1510), .S0(n1530) );
  HS65_GSS_XNOR2X3 U1598 ( .A(n1530), .B(n1515), .Z(\mul_b0/fa1_s0[6] ) );
  HS65_GS_AND2X4 U1599 ( .A(n1516), .B(n1891), .Z(\mul_b0/fa1_c0[20] ) );
  HS65_GS_AND2X4 U1600 ( .A(n1517), .B(x_z1[15]), .Z(\mul_b0/fa1_c0[19] ) );
  HS65_GS_AND2X4 U1601 ( .A(n1518), .B(n1891), .Z(\mul_b0/fa1_c0[18] ) );
  HS65_GS_AND2X4 U1602 ( .A(n1519), .B(x_z1[15]), .Z(\mul_b0/fa1_c0[17] ) );
  HS65_GS_AND2X4 U1603 ( .A(n1520), .B(n1891), .Z(\mul_b0/fa1_c0[16] ) );
  HS65_GS_AND2X4 U1604 ( .A(n1521), .B(x_z1[15]), .Z(\mul_b0/fa1_c0[15] ) );
  HS65_GS_AND2X4 U1605 ( .A(n1522), .B(x_z1[14]), .Z(\mul_b0/fa1_c0[14] ) );
  HS65_GS_AND2X4 U1606 ( .A(n1523), .B(x_z1[13]), .Z(\mul_b0/fa1_c0[13] ) );
  HS65_GS_AND2X4 U1607 ( .A(n1524), .B(x_z1[12]), .Z(\mul_b0/fa1_c0[12] ) );
  HS65_GS_AND2X4 U1608 ( .A(n1525), .B(x_z1[11]), .Z(\mul_b0/fa1_c0[11] ) );
  HS65_GS_AND2X4 U1609 ( .A(n1526), .B(x_z1[10]), .Z(\mul_b0/fa1_c0[10] ) );
  HS65_GS_AND2X4 U1610 ( .A(x_z1[9]), .B(n1527), .Z(\mul_b0/fa1_c0[9] ) );
  HS65_GS_AND2X4 U1611 ( .A(x_z1[8]), .B(n1528), .Z(\mul_b0/fa1_c0[8] ) );
  HS65_GS_AND2X4 U1612 ( .A(n1529), .B(x_z1[7]), .Z(\mul_b0/fa1_c0[7] ) );
  HS65_GS_AND2X4 U1613 ( .A(x_z1[6]), .B(n1530), .Z(\mul_b0/fa1_c0[6] ) );
  HS65_GS_AND2X4 U1614 ( .A(x_z1[5]), .B(x_z1[0]), .Z(\mul_b0/fa1_c0[5] ) );
  HS65_GS_FA1X4 U1615 ( .A0(n1533), .B0(n1532), .CI(n1531), .CO(n1029), .S0(
        n1534) );
  HS65_GS_AO12X4 U1616 ( .A(n1534), .B(n1554), .C(n1557), .Z(
        \mul_b0/result_sat[14] ) );
  HS65_GS_FA1X4 U1617 ( .A0(n1537), .B0(n1536), .CI(n1535), .CO(n1050), .S0(
        n1538) );
  HS65_GS_AO12X4 U1618 ( .A(n1538), .B(n1554), .C(n1557), .Z(
        \mul_b0/result_sat[10] ) );
  HS65_GS_FA1X4 U1619 ( .A0(n1541), .B0(n1540), .CI(n1539), .CO(n1537), .S0(
        n1542) );
  HS65_GS_AO12X4 U1620 ( .A(n1542), .B(n1554), .C(n1557), .Z(
        \mul_b0/result_sat[9] ) );
  HS65_GS_FA1X4 U1621 ( .A0(n1545), .B0(n1544), .CI(n1543), .CO(n1541), .S0(
        n1546) );
  HS65_GS_AO12X4 U1622 ( .A(n1546), .B(n1554), .C(n1557), .Z(
        \mul_b0/result_sat[8] ) );
  HS65_GS_FA1X4 U1623 ( .A0(n1549), .B0(n1548), .CI(n1547), .CO(n1545), .S0(
        n1550) );
  HS65_GS_AO12X4 U1624 ( .A(n1550), .B(n1554), .C(n1557), .Z(
        \mul_b0/result_sat[7] ) );
  HS65_GS_FA1X4 U1625 ( .A0(n1553), .B0(n1552), .CI(n1551), .CO(n1547), .S0(
        n1555) );
  HS65_GS_OA12X4 U1626 ( .A(n1557), .B(n1555), .C(n1554), .Z(
        \mul_b0/result_sat[6] ) );
  HS65_GS_AOI12X2 U1627 ( .A(n1560), .B(n1559), .C(n1556), .Z(n1558) );
  HS65_GS_CB4I6X4 U1628 ( .A(n1560), .B(n1559), .C(n1558), .D(n1557), .Z(
        \mul_b0/result_sat[5] ) );
  HS65_GS_OAI21X2 U1629 ( .A(n1562), .B(n1561), .C(n1579), .Z(n1563) );
  HS65_GS_OAI21X2 U1630 ( .A(n1565), .B(n1563), .C(n1868), .Z(
        \mul_a1/result_sat[1] ) );
  HS65_GS_FA1X4 U1631 ( .A0(n1566), .B0(n1565), .CI(n1564), .CO(n651), .S0(
        n1567) );
  HS65_GS_OA12X4 U1632 ( .A(n1581), .B(n1567), .C(n1579), .Z(
        \mul_a1/result_sat[2] ) );
  HS65_GS_FA1X4 U1633 ( .A0(n1570), .B0(n1569), .CI(n1568), .CO(n1573), .S0(
        n1571) );
  HS65_GS_OA12X4 U1634 ( .A(n1581), .B(n1571), .C(n1579), .Z(
        \mul_a1/result_sat[12] ) );
  HS65_GS_FA1X4 U1635 ( .A0(n1574), .B0(n1573), .CI(n1572), .CO(n1578), .S0(
        n1575) );
  HS65_GS_OA12X4 U1636 ( .A(n1581), .B(n1575), .C(n1579), .Z(
        \mul_a1/result_sat[13] ) );
  HS65_GS_FA1X4 U1637 ( .A0(n1578), .B0(n1577), .CI(n1576), .CO(n1074), .S0(
        n1580) );
  HS65_GS_OA12X4 U1638 ( .A(n1581), .B(n1580), .C(n1579), .Z(
        \mul_a1/result_sat[14] ) );
  HS65_GSS_XNOR2X3 U1639 ( .A(y_z1[0]), .B(n1843), .Z(\mul_a1/fa1_s2[14] ) );
  HS65_GSS_XNOR2X3 U1640 ( .A(n1628), .B(n1841), .Z(\mul_a1/fa1_s2[15] ) );
  HS65_GS_HA1X4 U1641 ( .A0(n1843), .B0(n1842), .CO(n1582), .S0(n1628) );
  HS65_GSS_XNOR2X3 U1642 ( .A(n1629), .B(n1839), .Z(\mul_a1/fa1_s2[16] ) );
  HS65_GS_HA1X4 U1643 ( .A0(n1841), .B0(n1582), .CO(n1583), .S0(n1629) );
  HS65_GSS_XNOR2X3 U1644 ( .A(n1630), .B(n1837), .Z(\mul_a1/fa1_s2[17] ) );
  HS65_GS_HA1X4 U1645 ( .A0(n1839), .B0(n1583), .CO(n1584), .S0(n1630) );
  HS65_GSS_XNOR2X3 U1646 ( .A(n1631), .B(n1835), .Z(\mul_a1/fa1_s2[18] ) );
  HS65_GS_HA1X4 U1647 ( .A0(n1837), .B0(n1584), .CO(n1585), .S0(n1631) );
  HS65_GSS_XNOR2X3 U1648 ( .A(n1632), .B(n1833), .Z(\mul_a1/fa1_s2[19] ) );
  HS65_GS_HA1X4 U1649 ( .A0(n1835), .B0(n1585), .CO(n1586), .S0(n1632) );
  HS65_GSS_XNOR2X3 U1650 ( .A(n1633), .B(n1831), .Z(\mul_a1/fa1_s2[20] ) );
  HS65_GS_HA1X4 U1651 ( .A0(n1833), .B0(n1586), .CO(n1587), .S0(n1633) );
  HS65_GSS_XNOR2X3 U1652 ( .A(n1634), .B(n1829), .Z(\mul_a1/fa1_s2[21] ) );
  HS65_GS_HA1X4 U1653 ( .A0(n1831), .B0(n1587), .CO(n1588), .S0(n1634) );
  HS65_GSS_XNOR2X3 U1654 ( .A(n1635), .B(n1827), .Z(\mul_a1/fa1_s2[22] ) );
  HS65_GS_HA1X4 U1655 ( .A0(n1829), .B0(n1588), .CO(n1589), .S0(n1635) );
  HS65_GSS_XNOR2X3 U1656 ( .A(n1636), .B(n1825), .Z(\mul_a1/fa1_s2[23] ) );
  HS65_GS_HA1X4 U1657 ( .A0(n1827), .B0(n1589), .CO(n1590), .S0(n1636) );
  HS65_GSS_XNOR2X3 U1658 ( .A(n1637), .B(n1823), .Z(\mul_a1/fa1_s2[24] ) );
  HS65_GS_HA1X4 U1659 ( .A0(n1825), .B0(n1590), .CO(n1591), .S0(n1637) );
  HS65_GSS_XNOR2X3 U1660 ( .A(n1797), .B(n1821), .Z(\mul_a1/fa1_s2[25] ) );
  HS65_GS_HA1X4 U1661 ( .A0(n1823), .B0(n1591), .CO(n1592), .S0(n1797) );
  HS65_GSS_XNOR2X3 U1662 ( .A(n1638), .B(n1819), .Z(\mul_a1/fa1_s2[26] ) );
  HS65_GS_HA1X4 U1663 ( .A0(n1821), .B0(n1592), .CO(n1593), .S0(n1638) );
  HS65_GSS_XNOR2X3 U1664 ( .A(n1639), .B(n1817), .Z(\mul_a1/fa1_s2[27] ) );
  HS65_GS_HA1X4 U1665 ( .A0(n1819), .B0(n1593), .CO(n1594), .S0(n1639) );
  HS65_GSS_XNOR2X3 U1666 ( .A(n1640), .B(n1815), .Z(\mul_a1/fa1_s2[28] ) );
  HS65_GS_HA1X4 U1667 ( .A0(n1817), .B0(n1594), .CO(n1595), .S0(n1640) );
  HS65_GSS_XNOR2X3 U1668 ( .A(n1641), .B(n1815), .Z(\mul_a1/fa1_s2[29] ) );
  HS65_GS_HA1X4 U1669 ( .A0(n1815), .B0(n1595), .CO(n1597), .S0(n1641) );
  HS65_GSS_XNOR2X3 U1670 ( .A(y_z1[15]), .B(n1597), .Z(n1596) );
  HS65_GSS_XNOR2X3 U1671 ( .A(n1596), .B(n1815), .Z(\mul_a1/fa1_s2[30] ) );
  HS65_GS_NOR2X2 U1672 ( .A(y_z1[15]), .B(n1597), .Z(n1598) );
  HS65_GSS_XNOR2X3 U1673 ( .A(n1598), .B(n1815), .Z(\mul_a1/fa1_s2[31] ) );
  HS65_GS_AND2X4 U1674 ( .A(y_z1[0]), .B(y_z1[3]), .Z(\mul_a1/fa1_c0[5] ) );
  HS65_GS_HA1X4 U1675 ( .A0(n1843), .B0(n1842), .CO(n1599), .S0(n1613) );
  HS65_GS_AND2X4 U1676 ( .A(n1613), .B(y_z1[4]), .Z(\mul_a1/fa1_c0[6] ) );
  HS65_GS_HA1X4 U1677 ( .A0(n1841), .B0(n1599), .CO(n1600), .S0(n1614) );
  HS65_GS_AND2X4 U1678 ( .A(n1614), .B(y_z1[5]), .Z(\mul_a1/fa1_c0[7] ) );
  HS65_GS_HA1X4 U1679 ( .A0(n1839), .B0(n1600), .CO(n1601), .S0(n1615) );
  HS65_GS_AND2X4 U1680 ( .A(n1615), .B(y_z1[6]), .Z(\mul_a1/fa1_c0[8] ) );
  HS65_GS_HA1X4 U1681 ( .A0(n1837), .B0(n1601), .CO(n1602), .S0(n1616) );
  HS65_GS_AND2X4 U1682 ( .A(n1616), .B(y_z1[7]), .Z(\mul_a1/fa1_c0[9] ) );
  HS65_GS_HA1X4 U1683 ( .A0(n1835), .B0(n1602), .CO(n1603), .S0(n1617) );
  HS65_GS_AND2X4 U1684 ( .A(n1617), .B(y_z1[8]), .Z(\mul_a1/fa1_c0[10] ) );
  HS65_GS_HA1X4 U1685 ( .A0(n1833), .B0(n1603), .CO(n1604), .S0(n1618) );
  HS65_GS_AND2X4 U1686 ( .A(n1618), .B(y_z1[9]), .Z(\mul_a1/fa1_c0[11] ) );
  HS65_GS_HA1X4 U1687 ( .A0(n1831), .B0(n1604), .CO(n1605), .S0(n1619) );
  HS65_GS_AND2X4 U1688 ( .A(n1619), .B(y_z1[10]), .Z(\mul_a1/fa1_c0[12] ) );
  HS65_GS_HA1X4 U1689 ( .A0(n1829), .B0(n1605), .CO(n1606), .S0(n1620) );
  HS65_GS_AND2X4 U1690 ( .A(n1620), .B(y_z1[11]), .Z(\mul_a1/fa1_c0[13] ) );
  HS65_GS_HA1X4 U1691 ( .A0(n1827), .B0(n1606), .CO(n1607), .S0(n1621) );
  HS65_GS_AND2X4 U1692 ( .A(n1621), .B(y_z1[12]), .Z(\mul_a1/fa1_c0[14] ) );
  HS65_GS_HA1X4 U1693 ( .A0(n1825), .B0(n1607), .CO(n1608), .S0(n1622) );
  HS65_GS_AND2X4 U1694 ( .A(n1622), .B(y_z1[13]), .Z(\mul_a1/fa1_c0[15] ) );
  HS65_GS_HA1X4 U1695 ( .A0(n1823), .B0(n1608), .CO(n1609), .S0(n1623) );
  HS65_GS_AND2X4 U1696 ( .A(n1623), .B(y_z1[14]), .Z(\mul_a1/fa1_c0[16] ) );
  HS65_GS_HA1X4 U1697 ( .A0(n1821), .B0(n1609), .CO(n1610), .S0(n1624) );
  HS65_GS_AND2X4 U1698 ( .A(n1624), .B(y_z1[15]), .Z(\mul_a1/fa1_c0[17] ) );
  HS65_GS_HA1X4 U1699 ( .A0(n1819), .B0(n1610), .CO(n1611), .S0(n1625) );
  HS65_GS_AND2X4 U1700 ( .A(n1625), .B(y_z1[15]), .Z(\mul_a1/fa1_c0[18] ) );
  HS65_GS_HA1X4 U1701 ( .A0(n1817), .B0(n1611), .CO(n1612), .S0(n1626) );
  HS65_GS_AND2X4 U1702 ( .A(n1626), .B(y_z1[15]), .Z(\mul_a1/fa1_c0[19] ) );
  HS65_GSS_XNOR2X3 U1703 ( .A(y_z1[15]), .B(n1612), .Z(n1627) );
  HS65_GS_AND2X4 U1704 ( .A(n1627), .B(y_z1[15]), .Z(\mul_a1/fa1_c0[20] ) );
  HS65_GSS_XNOR2X3 U1705 ( .A(n1613), .B(n1837), .Z(\mul_a1/fa1_s0[6] ) );
  HS65_GSS_XNOR2X3 U1706 ( .A(n1614), .B(n1835), .Z(\mul_a1/fa1_s0[7] ) );
  HS65_GSS_XNOR2X3 U1707 ( .A(n1615), .B(n1833), .Z(\mul_a1/fa1_s0[8] ) );
  HS65_GSS_XNOR2X3 U1708 ( .A(n1616), .B(n1831), .Z(\mul_a1/fa1_s0[9] ) );
  HS65_GSS_XNOR2X3 U1709 ( .A(n1617), .B(n1829), .Z(\mul_a1/fa1_s0[10] ) );
  HS65_GSS_XNOR2X3 U1710 ( .A(n1618), .B(n1827), .Z(\mul_a1/fa1_s0[11] ) );
  HS65_GSS_XNOR2X3 U1711 ( .A(n1619), .B(n1825), .Z(\mul_a1/fa1_s0[12] ) );
  HS65_GSS_XNOR2X3 U1712 ( .A(n1620), .B(n1823), .Z(\mul_a1/fa1_s0[13] ) );
  HS65_GSS_XNOR2X3 U1713 ( .A(n1621), .B(n1821), .Z(\mul_a1/fa1_s0[14] ) );
  HS65_GSS_XNOR2X3 U1714 ( .A(n1622), .B(n1819), .Z(\mul_a1/fa1_s0[15] ) );
  HS65_GSS_XNOR2X3 U1715 ( .A(n1623), .B(n1817), .Z(\mul_a1/fa1_s0[16] ) );
  HS65_GSS_XNOR2X3 U1716 ( .A(n1624), .B(n1815), .Z(\mul_a1/fa1_s0[17] ) );
  HS65_GSS_XNOR2X3 U1717 ( .A(n1625), .B(n1815), .Z(\mul_a1/fa1_s0[18] ) );
  HS65_GSS_XNOR2X3 U1718 ( .A(n1626), .B(n1815), .Z(\mul_a1/fa1_s0[19] ) );
  HS65_GSS_XNOR2X3 U1719 ( .A(n1627), .B(n1815), .Z(\mul_a1/fa1_s0[20] ) );
  HS65_GS_AND2X4 U1720 ( .A(y_z1[0]), .B(y_z1[1]), .Z(\mul_a1/fa1_c2[14] ) );
  HS65_GS_AND2X4 U1721 ( .A(n1628), .B(y_z1[2]), .Z(\mul_a1/fa1_c2[15] ) );
  HS65_GS_AND2X4 U1722 ( .A(n1629), .B(y_z1[3]), .Z(\mul_a1/fa1_c2[16] ) );
  HS65_GS_AND2X4 U1723 ( .A(n1630), .B(y_z1[4]), .Z(\mul_a1/fa1_c2[17] ) );
  HS65_GS_AND2X4 U1724 ( .A(n1631), .B(y_z1[5]), .Z(\mul_a1/fa1_c2[18] ) );
  HS65_GS_AND2X4 U1725 ( .A(n1632), .B(y_z1[6]), .Z(\mul_a1/fa1_c2[19] ) );
  HS65_GS_AND2X4 U1726 ( .A(n1633), .B(y_z1[7]), .Z(\mul_a1/fa1_c2[20] ) );
  HS65_GS_AND2X4 U1727 ( .A(n1634), .B(y_z1[8]), .Z(\mul_a1/fa1_c2[21] ) );
  HS65_GS_AND2X4 U1728 ( .A(n1635), .B(y_z1[9]), .Z(\mul_a1/fa1_c2[22] ) );
  HS65_GS_AND2X4 U1729 ( .A(n1636), .B(y_z1[10]), .Z(\mul_a1/fa1_c2[23] ) );
  HS65_GS_AND2X4 U1730 ( .A(n1637), .B(y_z1[11]), .Z(\mul_a1/fa1_c2[24] ) );
  HS65_GS_AND2X4 U1731 ( .A(n1638), .B(y_z1[13]), .Z(\mul_a1/fa1_c2[26] ) );
  HS65_GS_AND2X4 U1732 ( .A(n1639), .B(y_z1[14]), .Z(\mul_a1/fa1_c2[27] ) );
  HS65_GS_AND2X4 U1733 ( .A(n1640), .B(y_z1[15]), .Z(\mul_a1/fa1_c2[28] ) );
  HS65_GS_AND2X4 U1734 ( .A(n1641), .B(y_z1[15]), .Z(\mul_a1/fa1_c2[29] ) );
  HS65_GS_FA1X4 U1735 ( .A0(n1644), .B0(n1643), .CI(n1642), .CO(n1647), .S0(
        n1645) );
  HS65_GS_AO12X4 U1736 ( .A(n1645), .B(n1697), .C(n1699), .Z(
        \mul_a2/result_sat[1] ) );
  HS65_GS_FA1X4 U1737 ( .A0(n1648), .B0(n1647), .CI(n1646), .CO(n1651), .S0(
        n1649) );
  HS65_GS_OA12X4 U1738 ( .A(n1699), .B(n1649), .C(n1697), .Z(
        \mul_a2/result_sat[2] ) );
  HS65_GS_FA1X4 U1739 ( .A0(n1652), .B0(n1651), .CI(n1650), .CO(n1655), .S0(
        n1653) );
  HS65_GS_AO12X4 U1740 ( .A(n1653), .B(n1697), .C(n1699), .Z(
        \mul_a2/result_sat[3] ) );
  HS65_GS_FA1X4 U1741 ( .A0(n1656), .B0(n1655), .CI(n1654), .CO(n1659), .S0(
        n1657) );
  HS65_GS_AO12X4 U1742 ( .A(n1657), .B(n1697), .C(n1699), .Z(
        \mul_a2/result_sat[4] ) );
  HS65_GS_FA1X4 U1743 ( .A0(n1660), .B0(n1659), .CI(n1658), .CO(n1663), .S0(
        n1661) );
  HS65_GS_OA12X4 U1744 ( .A(n1699), .B(n1661), .C(n1697), .Z(
        \mul_a2/result_sat[5] ) );
  HS65_GS_FA1X4 U1745 ( .A0(n1664), .B0(n1663), .CI(n1662), .CO(n1667), .S0(
        n1665) );
  HS65_GS_AO12X4 U1746 ( .A(n1665), .B(n1697), .C(n1699), .Z(
        \mul_a2/result_sat[6] ) );
  HS65_GS_FA1X4 U1747 ( .A0(n1668), .B0(n1667), .CI(n1666), .CO(n1671), .S0(
        n1669) );
  HS65_GS_OA12X4 U1748 ( .A(n1699), .B(n1669), .C(n1697), .Z(
        \mul_a2/result_sat[7] ) );
  HS65_GS_FA1X4 U1749 ( .A0(n1672), .B0(n1671), .CI(n1670), .CO(n1675), .S0(
        n1673) );
  HS65_GS_AO12X4 U1750 ( .A(n1673), .B(n1697), .C(n1699), .Z(
        \mul_a2/result_sat[8] ) );
  HS65_GS_FA1X4 U1751 ( .A0(n1676), .B0(n1675), .CI(n1674), .CO(n1680), .S0(
        n1677) );
  HS65_GS_OA12X4 U1752 ( .A(n1699), .B(n1677), .C(n1697), .Z(
        \mul_a2/result_sat[9] ) );
  HS65_GS_FA1X4 U1753 ( .A0(n1680), .B0(n1679), .CI(n1678), .CO(n1683), .S0(
        n1681) );
  HS65_GS_OA12X4 U1754 ( .A(n1699), .B(n1681), .C(n1697), .Z(
        \mul_a2/result_sat[10] ) );
  HS65_GS_FA1X4 U1755 ( .A0(n1684), .B0(n1683), .CI(n1682), .CO(n1687), .S0(
        n1685) );
  HS65_GS_OA12X4 U1756 ( .A(n1699), .B(n1685), .C(n1697), .Z(
        \mul_a2/result_sat[11] ) );
  HS65_GS_FA1X4 U1757 ( .A0(n1688), .B0(n1687), .CI(n1686), .CO(n1691), .S0(
        n1689) );
  HS65_GS_OA12X4 U1758 ( .A(n1699), .B(n1689), .C(n1697), .Z(
        \mul_a2/result_sat[12] ) );
  HS65_GS_FA1X4 U1759 ( .A0(n1692), .B0(n1691), .CI(n1690), .CO(n1696), .S0(
        n1693) );
  HS65_GS_OA12X4 U1760 ( .A(n1699), .B(n1693), .C(n1697), .Z(
        \mul_a2/result_sat[13] ) );
  HS65_GS_FA1X4 U1761 ( .A0(n1696), .B0(n1695), .CI(n1694), .CO(n1121), .S0(
        n1698) );
  HS65_GS_OA12X4 U1762 ( .A(n1699), .B(n1698), .C(n1697), .Z(
        \mul_a2/result_sat[14] ) );
  HS65_GSS_XNOR2X3 U1763 ( .A(n1700), .B(n1314), .Z(\mul_a2/fa1_s2[14] ) );
  HS65_GSS_XNOR2X3 U1764 ( .A(n1701), .B(n1844), .Z(\mul_a2/fa1_s2[15] ) );
  HS65_GSS_XNOR2X3 U1765 ( .A(n1703), .B(n1702), .Z(\mul_a2/fa1_s2[16] ) );
  HS65_GSS_XNOR2X3 U1766 ( .A(n1705), .B(n1704), .Z(\mul_a2/fa1_s2[17] ) );
  HS65_GSS_XNOR2X3 U1767 ( .A(n1707), .B(n1706), .Z(\mul_a2/fa1_s2[18] ) );
  HS65_GSS_XNOR2X3 U1768 ( .A(n1709), .B(n1708), .Z(\mul_a2/fa1_s2[19] ) );
  HS65_GSS_XNOR2X3 U1769 ( .A(n1711), .B(n1710), .Z(\mul_a2/fa1_s2[20] ) );
  HS65_GSS_XNOR2X3 U1770 ( .A(n1713), .B(n1712), .Z(\mul_a2/fa1_s2[21] ) );
  HS65_GSS_XNOR2X3 U1771 ( .A(n1715), .B(n1714), .Z(\mul_a2/fa1_s2[22] ) );
  HS65_GSS_XNOR2X3 U1772 ( .A(n1717), .B(n1716), .Z(\mul_a2/fa1_s2[23] ) );
  HS65_GSS_XNOR2X3 U1773 ( .A(n1719), .B(n1718), .Z(\mul_a2/fa1_s2[24] ) );
  HS65_GSS_XNOR2X3 U1774 ( .A(n1721), .B(n1720), .Z(\mul_a2/fa1_s2[25] ) );
  HS65_GSS_XNOR2X3 U1775 ( .A(n1723), .B(n1722), .Z(\mul_a2/fa1_s2[26] ) );
  HS65_GSS_XNOR2X3 U1776 ( .A(n1725), .B(n1724), .Z(\mul_a2/fa1_s2[27] ) );
  HS65_GSS_XNOR2X3 U1777 ( .A(n1727), .B(n1726), .Z(\mul_a2/fa1_s2[28] ) );
  HS65_GS_AND2X4 U1778 ( .A(n1728), .B(\mul_a2/fa1_s0[0] ), .Z(
        \mul_a2/fa1_c1[8] ) );
  HS65_GS_AND2X4 U1779 ( .A(n1730), .B(n1729), .Z(\mul_a2/fa1_c1[9] ) );
  HS65_GS_PAO2X4 U1780 ( .A(n1732), .B(n1731), .P(\mul_a2/fa1_s0[0] ), .Z(
        \mul_a2/fa1_c1[10] ) );
  HS65_GS_PAO2X4 U1781 ( .A(n1734), .B(n1733), .P(\mul_a2/fa1_s0[1] ), .Z(
        \mul_a2/fa1_c1[11] ) );
  HS65_GS_PAO2X4 U1782 ( .A(n1736), .B(n1735), .P(y_z2[2]), .Z(
        \mul_a2/fa1_c1[12] ) );
  HS65_GS_HA1X4 U1783 ( .A0(n1738), .B0(n1737), .CO(n1762), .S0(n1761) );
  HS65_GS_AND2X4 U1784 ( .A(n1761), .B(x_z2[8]), .Z(\mul_b1/fa1_c0[8] ) );
  HS65_GS_HA1X4 U1785 ( .A0(n1756), .B0(n1739), .CO(n1740), .S0(n1766) );
  HS65_GS_AND2X4 U1786 ( .A(n1766), .B(x_z2[10]), .Z(\mul_b1/fa1_c0[10] ) );
  HS65_GS_HA1X4 U1787 ( .A0(n1758), .B0(n1740), .CO(n1743), .S0(n1768) );
  HS65_GS_AND2X4 U1788 ( .A(n1768), .B(x_z2[11]), .Z(\mul_b1/fa1_c0[11] ) );
  HS65_GS_HA1X4 U1789 ( .A0(n1742), .B0(n1741), .CO(n1737), .S0(n1759) );
  HS65_GS_AND2X4 U1790 ( .A(n1759), .B(x_z2[7]), .Z(\mul_b1/fa1_c0[7] ) );
  HS65_GS_HA1X4 U1791 ( .A0(n1760), .B0(n1743), .CO(n1744), .S0(n1770) );
  HS65_GS_AND2X4 U1792 ( .A(n1770), .B(x_z2[12]), .Z(\mul_b1/fa1_c0[12] ) );
  HS65_GS_HA1X4 U1793 ( .A0(n1764), .B0(n1744), .CO(n1745), .S0(n1772) );
  HS65_GS_AND2X4 U1794 ( .A(n1772), .B(x_z2[13]), .Z(\mul_b1/fa1_c0[13] ) );
  HS65_GS_HA1X4 U1795 ( .A0(n1765), .B0(n1745), .CO(n1748), .S0(n1774) );
  HS65_GS_AND2X4 U1796 ( .A(n1774), .B(x_z2[14]), .Z(\mul_b1/fa1_c0[14] ) );
  HS65_GS_HA1X4 U1797 ( .A0(n1747), .B0(n1746), .CO(n1741), .S0(n1757) );
  HS65_GS_AND2X4 U1798 ( .A(n1757), .B(x_z2[6]), .Z(\mul_b1/fa1_c0[6] ) );
  HS65_GS_HA1X4 U1799 ( .A0(n1767), .B0(n1748), .CO(n1751), .S0(n1775) );
  HS65_GS_AND2X4 U1800 ( .A(n1775), .B(x_z2[15]), .Z(\mul_b1/fa1_c0[15] ) );
  HS65_GS_HA1X4 U1801 ( .A0(n1750), .B0(n1749), .CO(n1746), .S0(n1755) );
  HS65_GS_AND2X4 U1802 ( .A(n1755), .B(x_z2[5]), .Z(\mul_b1/fa1_c0[5] ) );
  HS65_GS_HA1X4 U1803 ( .A0(n1769), .B0(n1751), .CO(n1752), .S0(n1776) );
  HS65_GS_AND2X4 U1804 ( .A(n1776), .B(x_z2[15]), .Z(\mul_b1/fa1_c0[16] ) );
  HS65_GS_AND2X4 U1805 ( .A(x_z2[0]), .B(x_z2[4]), .Z(\mul_b1/fa1_c0[4] ) );
  HS65_GS_HA1X4 U1806 ( .A0(n1771), .B0(n1752), .CO(n1753), .S0(n1777) );
  HS65_GS_AND2X4 U1807 ( .A(n1777), .B(x_z2[15]), .Z(\mul_b1/fa1_c0[17] ) );
  HS65_GS_HA1X4 U1808 ( .A0(n1773), .B0(n1753), .CO(n1754), .S0(n1778) );
  HS65_GS_AND2X4 U1809 ( .A(n1778), .B(x_z2[15]), .Z(\mul_b1/fa1_c0[18] ) );
  HS65_GS_HA1X4 U1810 ( .A0(n1810), .B0(n1754), .CO(n1780), .S0(n1779) );
  HS65_GS_AND2X4 U1811 ( .A(n1779), .B(x_z2[15]), .Z(\mul_b1/fa1_c0[19] ) );
  HS65_GSS_XNOR2X3 U1812 ( .A(n1755), .B(n1763), .Z(\mul_b1/fa1_s0[5] ) );
  HS65_GSS_XNOR2X3 U1813 ( .A(n1757), .B(n1756), .Z(\mul_b1/fa1_s0[6] ) );
  HS65_GSS_XNOR2X3 U1814 ( .A(n1759), .B(n1758), .Z(\mul_b1/fa1_s0[7] ) );
  HS65_GSS_XNOR2X3 U1815 ( .A(n1761), .B(n1760), .Z(\mul_b1/fa1_s0[8] ) );
  HS65_GS_HA1X4 U1816 ( .A0(n1763), .B0(n1762), .CO(n1739), .S0(n1798) );
  HS65_GSS_XNOR2X3 U1817 ( .A(n1798), .B(n1764), .Z(\mul_b1/fa1_s0[9] ) );
  HS65_GSS_XNOR2X3 U1818 ( .A(n1766), .B(n1765), .Z(\mul_b1/fa1_s0[10] ) );
  HS65_GSS_XNOR2X3 U1819 ( .A(n1768), .B(n1767), .Z(\mul_b1/fa1_s0[11] ) );
  HS65_GSS_XNOR2X3 U1820 ( .A(n1770), .B(n1769), .Z(\mul_b1/fa1_s0[12] ) );
  HS65_GSS_XNOR2X3 U1821 ( .A(n1772), .B(n1771), .Z(\mul_b1/fa1_s0[13] ) );
  HS65_GSS_XNOR2X3 U1822 ( .A(n1774), .B(n1773), .Z(\mul_b1/fa1_s0[14] ) );
  HS65_GSS_XNOR2X3 U1823 ( .A(n1775), .B(n1810), .Z(\mul_b1/fa1_s0[15] ) );
  HS65_GSS_XNOR2X3 U1824 ( .A(n1776), .B(n1810), .Z(\mul_b1/fa1_s0[16] ) );
  HS65_GSS_XNOR2X3 U1825 ( .A(n1777), .B(n1810), .Z(\mul_b1/fa1_s0[17] ) );
  HS65_GSS_XNOR2X3 U1826 ( .A(n1778), .B(n1810), .Z(\mul_b1/fa1_s0[18] ) );
  HS65_GSS_XNOR2X3 U1827 ( .A(n1779), .B(n1810), .Z(\mul_b1/fa1_s0[19] ) );
  HS65_GSS_XNOR2X3 U1828 ( .A(x_z2[15]), .B(n1780), .Z(n1781) );
  HS65_GSS_XNOR2X3 U1829 ( .A(n1781), .B(n1810), .Z(\mul_b1/fa1_s0[20] ) );
  HS65_GS_AND2X4 U1830 ( .A(n1782), .B(x_z2[0]), .Z(\mul_b1/fa1_c2[14] ) );
  HS65_GS_AND2X4 U1831 ( .A(n1783), .B(x_z2[1]), .Z(\mul_b1/fa1_c2[15] ) );
  HS65_GS_AND2X4 U1832 ( .A(n1784), .B(x_z2[2]), .Z(\mul_b1/fa1_c2[16] ) );
  HS65_GS_AND2X4 U1833 ( .A(n1785), .B(x_z2[3]), .Z(\mul_b1/fa1_c2[17] ) );
  HS65_GS_AND2X4 U1834 ( .A(n1786), .B(x_z2[4]), .Z(\mul_b1/fa1_c2[18] ) );
  HS65_GS_AND2X4 U1835 ( .A(n1787), .B(x_z2[5]), .Z(\mul_b1/fa1_c2[19] ) );
  HS65_GS_AND2X4 U1836 ( .A(n1788), .B(x_z2[6]), .Z(\mul_b1/fa1_c2[20] ) );
  HS65_GS_AND2X4 U1837 ( .A(n1789), .B(x_z2[7]), .Z(\mul_b1/fa1_c2[21] ) );
  HS65_GS_AND2X4 U1838 ( .A(n1790), .B(x_z2[8]), .Z(\mul_b1/fa1_c2[22] ) );
  HS65_GS_AND2X4 U1839 ( .A(n1791), .B(x_z2[9]), .Z(\mul_b1/fa1_c2[23] ) );
  HS65_GS_AND2X4 U1840 ( .A(n1792), .B(x_z2[10]), .Z(\mul_b1/fa1_c2[24] ) );
  HS65_GS_AND2X4 U1841 ( .A(n1793), .B(x_z2[11]), .Z(\mul_b1/fa1_c2[25] ) );
  HS65_GS_AND2X4 U1842 ( .A(n1794), .B(x_z2[12]), .Z(\mul_b1/fa1_c2[26] ) );
  HS65_GS_AND2X4 U1843 ( .A(n1795), .B(x_z2[13]), .Z(\mul_b1/fa1_c2[27] ) );
  HS65_GS_AND2X4 U1844 ( .A(n1796), .B(x_z2[14]), .Z(\mul_b1/fa1_c2[28] ) );
  HS65_GS_AND2X4 U1845 ( .A(n1797), .B(y_z1[12]), .Z(\mul_a1/fa1_c2[25] ) );
  HS65_GS_AND2X4 U1846 ( .A(n1798), .B(x_z2[9]), .Z(\mul_b1/fa1_c0[9] ) );
  HS65_GS_AOI12X2 U1847 ( .A(n1802), .B(n1801), .C(n1799), .Z(n1800) );
  HS65_GS_CB4I6X4 U1848 ( .A(n1802), .B(n1801), .C(n1800), .D(n1806), .Z(
        \mul_b2/result_sat[13] ) );
  HS65_GS_FA1X4 U1849 ( .A0(n1805), .B0(n1804), .CI(n1803), .CO(n1151), .S0(
        n1808) );
  HS65_GS_AO12X4 U1850 ( .A(n1808), .B(n1807), .C(n1806), .Z(
        \mul_b2/result_sat[14] ) );
  HS65_GS_NOR2X2 U1851 ( .A(x_z2[15]), .B(n1809), .Z(n1811) );
  HS65_GSS_XNOR2X3 U1852 ( .A(n1811), .B(n1810), .Z(\mul_b1/fa1_s2[29] ) );
  HS65_GS_AND2X4 U1853 ( .A(\mul_a2/fa1_s0[0] ), .B(y_z2[2]), .Z(n1885) );
  HS65_GS_AND2X4 U1854 ( .A(n1812), .B(y_z2[3]), .Z(n1887) );
  HS65_GSS_XNOR2X3 U1855 ( .A(y_z1[15]), .B(n1813), .Z(\C53/DATA4_24 ) );
  HS65_GS_HA1X4 U1856 ( .A0(n1815), .B0(n1814), .CO(n1813), .S0(\C53/DATA4_23 ) );
  HS65_GS_HA1X4 U1857 ( .A0(n1817), .B0(n1816), .CO(n1814), .S0(\C53/DATA4_22 ) );
  HS65_GS_HA1X4 U1858 ( .A0(n1819), .B0(n1818), .CO(n1816), .S0(\C53/DATA4_21 ) );
  HS65_GS_HA1X4 U1859 ( .A0(n1821), .B0(n1820), .CO(n1818), .S0(\C53/DATA4_20 ) );
  HS65_GS_HA1X4 U1860 ( .A0(n1823), .B0(n1822), .CO(n1820), .S0(\C53/DATA4_19 ) );
  HS65_GS_HA1X4 U1861 ( .A0(n1825), .B0(n1824), .CO(n1822), .S0(\C53/DATA4_18 ) );
  HS65_GS_HA1X4 U1862 ( .A0(n1827), .B0(n1826), .CO(n1824), .S0(\C53/DATA4_17 ) );
  HS65_GS_HA1X4 U1863 ( .A0(n1829), .B0(n1828), .CO(n1826), .S0(\C53/DATA4_16 ) );
  HS65_GS_HA1X4 U1864 ( .A0(n1831), .B0(n1830), .CO(n1828), .S0(\C53/DATA4_15 ) );
  HS65_GS_HA1X4 U1865 ( .A0(n1833), .B0(n1832), .CO(n1830), .S0(\C53/DATA4_14 ) );
  HS65_GS_HA1X4 U1866 ( .A0(n1835), .B0(n1834), .CO(n1832), .S0(\C53/DATA4_13 ) );
  HS65_GS_HA1X4 U1867 ( .A0(n1837), .B0(n1836), .CO(n1834), .S0(\C53/DATA4_12 ) );
  HS65_GS_HA1X4 U1868 ( .A0(n1839), .B0(n1838), .CO(n1836), .S0(\C53/DATA4_11 ) );
  HS65_GS_HA1X4 U1869 ( .A0(n1841), .B0(n1840), .CO(n1838), .S0(\C53/DATA4_10 ) );
  HS65_GS_HA1X4 U1870 ( .A0(n1843), .B0(n1842), .CO(n1840), .S0(\C53/DATA4_9 )
         );
  HS65_GS_HA1X4 U1871 ( .A0(n1844), .B0(n1314), .CO(n1315), .S0(
        \mul_a2/fa1_s1[7] ) );
  HS65_GS_PAOI2X1 U1872 ( .A(n1850), .B(n1848), .P(n1847), .Z(
        \mul_b2/fa1_c0[4] ) );
  HS65_GS_PAOI2X1 U1873 ( .A(n1851), .B(n1846), .P(n1845), .Z(
        \mul_b2/fa1_c0[5] ) );
  HS65_GS_AOI12X2 U1874 ( .A(n1848), .B(n1847), .C(\mul_b2/fa1_c0[2] ), .Z(
        n1849) );
  HS65_GS_MUXI21X2 U1875 ( .D0(n1850), .D1(x_reg2[4]), .S0(n1849), .Z(
        \mul_b2/fa1_s0[4] ) );
  HS65_GS_MUXI21X2 U1876 ( .D0(n1851), .D1(x_reg2[5]), .S0(\mul_b2/fa1_s0[3] ), 
        .Z(\mul_b2/fa1_s0[5] ) );
  HS65_GS_FA1X4 U1877 ( .A0(x_reg2[6]), .B0(x_reg2[4]), .CI(x_reg2[2]), .CO(
        \mul_b2/fa1_c0[6] ), .S0(\mul_b2/fa1_s0[6] ) );
  HS65_GS_FA1X4 U1878 ( .A0(x_reg2[7]), .B0(x_reg2[5]), .CI(x_reg2[3]), .CO(
        \mul_b2/fa1_c0[7] ), .S0(\mul_b2/fa1_s0[7] ) );
  HS65_GS_FA1X4 U1879 ( .A0(x_reg2[8]), .B0(x_reg2[6]), .CI(x_reg2[4]), .CO(
        \mul_b2/fa1_c0[8] ), .S0(\mul_b2/fa1_s0[8] ) );
  HS65_GS_FA1X4 U1880 ( .A0(x_reg2[9]), .B0(x_reg2[7]), .CI(x_reg2[5]), .CO(
        \mul_b2/fa1_c0[9] ), .S0(\mul_b2/fa1_s0[9] ) );
  HS65_GS_FA1X4 U1881 ( .A0(x_reg2[10]), .B0(x_reg2[8]), .CI(x_reg2[6]), .CO(
        \mul_b2/fa1_c0[10] ), .S0(\mul_b2/fa1_s0[10] ) );
  HS65_GS_FA1X4 U1882 ( .A0(x_reg2[11]), .B0(x_reg2[9]), .CI(x_reg2[7]), .CO(
        \mul_b2/fa1_c0[11] ), .S0(\mul_b2/fa1_s0[11] ) );
  HS65_GS_FA1X4 U1883 ( .A0(x_reg2[12]), .B0(x_reg2[10]), .CI(x_reg2[8]), .CO(
        \mul_b2/fa1_c0[12] ), .S0(\mul_b2/fa1_s0[12] ) );
  HS65_GS_FA1X4 U1884 ( .A0(x_reg2[13]), .B0(x_reg2[11]), .CI(x_reg2[9]), .CO(
        \mul_b2/fa1_c0[13] ), .S0(\mul_b2/fa1_s0[13] ) );
  HS65_GS_FA1X4 U1885 ( .A0(x_reg2[14]), .B0(x_reg2[12]), .CI(x_reg2[10]), 
        .CO(\mul_b2/fa1_c0[14] ), .S0(\mul_b2/fa1_s0[14] ) );
  HS65_GS_FA1X4 U1886 ( .A0(n1889), .B0(x_reg2[13]), .CI(x_reg2[11]), .CO(
        \mul_b2/fa1_c0[15] ), .S0(\mul_b2/fa1_s0[15] ) );
  HS65_GS_FA1X4 U1887 ( .A0(n1889), .B0(x_reg2[14]), .CI(x_reg2[12]), .CO(
        \mul_b2/fa1_c0[16] ), .S0(\mul_b2/fa1_s0[16] ) );
  HS65_GS_FA1X4 U1888 ( .A0(n1854), .B0(n1853), .CI(n1852), .CO(n1856), .S0(
        n1855) );
  HS65_GS_AOI12X2 U1889 ( .A(n1855), .B(n1868), .C(n1867), .Z(
        \mul_a1/result_sat[6] ) );
  HS65_GS_FA1X4 U1890 ( .A0(n1858), .B0(n1857), .CI(n1856), .CO(n1109), .S0(
        n1859) );
  HS65_GS_AOI12X2 U1891 ( .A(n1859), .B(n1868), .C(n1867), .Z(
        \mul_a1/result_sat[7] ) );
  HS65_GS_AOI12X2 U1892 ( .A(n1862), .B(n1861), .C(n1860), .Z(n1863) );
  HS65_GS_AOI12X2 U1893 ( .A(n1863), .B(n1868), .C(n1867), .Z(
        \mul_a1/result_sat[9] ) );
  HS65_GS_AOI12X2 U1894 ( .A(n1866), .B(n1865), .C(n1864), .Z(n1869) );
  HS65_GS_AOI12X2 U1895 ( .A(n1869), .B(n1868), .C(n1867), .Z(
        \mul_a1/result_sat[10] ) );
  HS65_GS_CBI4I1X3 U1896 ( .A(n1872), .B(n1871), .C(n1870), .D(n1880), .Z(
        n1873) );
  HS65_GS_AND2X4 U1897 ( .A(n1873), .B(n1878), .Z(\mul_b1/result_sat[0] ) );
  HS65_GS_NOR2X2 U1898 ( .A(n1875), .B(n1874), .Z(n1876) );
  HS65_GSS_XNOR2X3 U1899 ( .A(n1877), .B(n1876), .Z(n1881) );
  HS65_GS_IVX2 U1900 ( .A(n1878), .Z(n1879) );
  HS65_GS_AOI12X2 U1901 ( .A(n1881), .B(n1880), .C(n1879), .Z(
        \mul_b1/result_sat[14] ) );
  HS65_GS_AOI12X2 U1902 ( .A(n1884), .B(n1883), .C(n1882), .Z(n1941) );
endmodule


module opti_sos_2 ( clk, rst_n, data_in, valid_in, b0, b1, b2, a1, a2, 
        data_out, valid_out );
  input [15:0] data_in;
  input [15:0] b0;
  input [15:0] b1;
  input [15:0] b2;
  input [15:0] a1;
  input [15:0] a2;
  output [15:0] data_out;
  input clk, rst_n, valid_in;
  output valid_out;
  wire   valid_T1, valid_T3, valid_T2, \mul_b0/result_sat[15] ,
         \mul_b0/result_sat[14] , \mul_b0/result_sat[13] ,
         \mul_b0/result_sat[12] , \mul_b0/result_sat[11] ,
         \mul_b0/result_sat[10] , \mul_b0/result_sat[9] ,
         \mul_b0/result_sat[8] , \mul_b0/result_sat[7] ,
         \mul_b0/result_sat[6] , \mul_b0/result_sat[5] ,
         \mul_b0/result_sat[4] , \mul_b0/result_sat[3] ,
         \mul_b0/result_sat[2] , \mul_b0/result_sat[1] ,
         \mul_b0/result_sat[0] , \mul_b0/fa1_s2_r[33] , \mul_b0/fa1_s2_r[32] ,
         \mul_b0/fa1_s2_r[31] , \mul_b0/fa1_s2_r[30] , \mul_b0/fa1_s2_r[29] ,
         \mul_b0/fa1_s2_r[28] , \mul_b0/fa1_s2_r[27] , \mul_b0/fa1_s2_r[26] ,
         \mul_b0/fa1_s2_r[25] , \mul_b0/fa1_s2_r[24] , \mul_b0/fa1_s2_r[23] ,
         \mul_b0/fa1_s2_r[22] , \mul_b0/fa1_s2_r[21] , \mul_b0/fa1_s2_r[20] ,
         \mul_b0/fa1_s2_r[19] , \mul_b0/fa1_s2_r[18] , \mul_b0/fa1_s2_r[17] ,
         \mul_b0/fa1_s2_r[16] , \mul_b0/fa1_s2_r[15] , \mul_b0/fa1_s2_r[14] ,
         \mul_b0/fa1_s2_r[13] , \mul_b0/fa1_s2_r[12] , \mul_b0/fa1_s1_r[33] ,
         \mul_b0/fa1_s1_r[32] , \mul_b0/fa1_s1_r[31] , \mul_b0/fa1_s1_r[30] ,
         \mul_b0/fa1_s1_r[29] , \mul_b0/fa1_s1_r[28] , \mul_b0/fa1_s1_r[27] ,
         \mul_b0/fa1_s1_r[26] , \mul_b0/fa1_s1_r[25] , \mul_b0/fa1_s1_r[24] ,
         \mul_b0/fa1_s1_r[23] , \mul_b0/fa1_s1_r[22] , \mul_b0/fa1_s1_r[21] ,
         \mul_b0/fa1_s1_r[20] , \mul_b0/fa1_s1_r[19] , \mul_b0/fa1_s1_r[18] ,
         \mul_b0/fa1_s1_r[17] , \mul_b0/fa1_s1_r[16] , \mul_b0/fa1_s1_r[15] ,
         \mul_b0/fa1_s1_r[14] , \mul_b0/fa1_s1_r[13] , \mul_b0/fa1_s1_r[12] ,
         \mul_b0/fa1_s1_r[11] , \mul_b0/fa1_s1_r[10] , \mul_b0/fa1_s1_r[9] ,
         \mul_b0/fa1_s1_r[8] , \mul_b0/fa1_c0_r[20] , \mul_b0/fa1_c0_r[19] ,
         \mul_b0/fa1_c0_r[18] , \mul_b0/fa1_c0_r[17] , \mul_b0/fa1_c0_r[16] ,
         \mul_b0/fa1_c0_r[15] , \mul_b0/fa1_c0_r[14] , \mul_b0/fa1_c0_r[13] ,
         \mul_b0/fa1_c0_r[12] , \mul_b0/fa1_c0_r[11] , \mul_b0/fa1_c0_r[10] ,
         \mul_b0/fa1_c0_r[9] , \mul_b0/fa1_c0_r[8] , \mul_b0/fa1_c0_r[7] ,
         \mul_b0/fa1_c0_r[6] , \mul_b0/fa1_c0_r[5] , \mul_b0/fa1_s0_r[33] ,
         \mul_b0/fa1_s0_r[32] , \mul_b0/fa1_s0_r[31] , \mul_b0/fa1_s0_r[30] ,
         \mul_b0/fa1_s0_r[29] , \mul_b0/fa1_s0_r[28] , \mul_b0/fa1_s0_r[27] ,
         \mul_b0/fa1_s0_r[26] , \mul_b0/fa1_s0_r[25] , \mul_b0/fa1_s0_r[24] ,
         \mul_b0/fa1_s0_r[23] , \mul_b0/fa1_s0_r[22] , \mul_b0/fa1_s0_r[21] ,
         \mul_b0/fa1_s0_r[20] , \mul_b0/fa1_s0_r[19] , \mul_b0/fa1_s0_r[18] ,
         \mul_b0/fa1_s0_r[17] , \mul_b0/fa1_s0_r[16] , \mul_b0/fa1_s0_r[15] ,
         \mul_b0/fa1_s0_r[14] , \mul_b0/fa1_s0_r[13] , \mul_b0/fa1_s0_r[12] ,
         \mul_b0/fa1_s0_r[11] , \mul_b0/fa1_s0_r[10] , \mul_b0/fa1_s0_r[9] ,
         \mul_b0/fa1_s0_r[8] , \mul_b0/fa1_s0_r[7] , \mul_b0/fa1_s0_r[6] ,
         \mul_b0/fa1_c0[20] , \mul_b0/fa1_c0[19] , \mul_b0/fa1_c0[18] ,
         \mul_b0/fa1_c0[17] , \mul_b0/fa1_c0[16] , \mul_b0/fa1_c0[15] ,
         \mul_b0/fa1_c0[14] , \mul_b0/fa1_c0[13] , \mul_b0/fa1_c0[12] ,
         \mul_b0/fa1_c0[11] , \mul_b0/fa1_c0[10] , \mul_b0/fa1_c0[9] ,
         \mul_b0/fa1_c0[8] , \mul_b0/fa1_c0[7] , \mul_b0/fa1_c0[6] ,
         \mul_b0/fa1_c0[5] , \mul_b0/fa1_s0[31] , \mul_b0/fa1_s0[20] ,
         \mul_b0/fa1_s0[19] , \mul_b0/fa1_s0[18] , \mul_b0/fa1_s0[17] ,
         \mul_b0/fa1_s0[16] , \mul_b0/fa1_s0[15] , \mul_b0/fa1_s0[14] ,
         \mul_b0/fa1_s0[13] , \mul_b0/fa1_s0[12] , \mul_b0/fa1_s0[11] ,
         \mul_b0/fa1_s0[10] , \mul_b0/fa1_s0[9] , \mul_b0/fa1_s0[8] ,
         \mul_b0/fa1_s0[7] , \mul_b0/fa1_s0[6] , \mul_b1/result_sat[15] ,
         \mul_b1/result_sat[14] , \mul_b1/result_sat[13] ,
         \mul_b1/result_sat[12] , \mul_b1/result_sat[11] ,
         \mul_b1/result_sat[10] , \mul_b1/result_sat[9] ,
         \mul_b1/result_sat[8] , \mul_b1/result_sat[7] ,
         \mul_b1/result_sat[6] , \mul_b1/result_sat[5] ,
         \mul_b1/result_sat[4] , \mul_b1/result_sat[3] ,
         \mul_b1/result_sat[2] , \mul_b1/result_sat[1] ,
         \mul_b1/result_sat[0] , \mul_b1/fa1_c2_r[28] , \mul_b1/fa1_c2_r[27] ,
         \mul_b1/fa1_c2_r[26] , \mul_b1/fa1_c2_r[25] , \mul_b1/fa1_c2_r[24] ,
         \mul_b1/fa1_c2_r[23] , \mul_b1/fa1_c2_r[22] , \mul_b1/fa1_c2_r[21] ,
         \mul_b1/fa1_c2_r[20] , \mul_b1/fa1_c2_r[19] , \mul_b1/fa1_c2_r[18] ,
         \mul_b1/fa1_c2_r[17] , \mul_b1/fa1_c2_r[16] , \mul_b1/fa1_c2_r[15] ,
         \mul_b1/fa1_c2_r[14] , \mul_b1/fa1_s2_r[33] , \mul_b1/fa1_s2_r[32] ,
         \mul_b1/fa1_s2_r[31] , \mul_b1/fa1_s2_r[30] , \mul_b1/fa1_s2_r[29] ,
         \mul_b1/fa1_s2_r[28] , \mul_b1/fa1_s2_r[27] , \mul_b1/fa1_s2_r[26] ,
         \mul_b1/fa1_s2_r[25] , \mul_b1/fa1_s2_r[24] , \mul_b1/fa1_s2_r[23] ,
         \mul_b1/fa1_s2_r[22] , \mul_b1/fa1_s2_r[21] , \mul_b1/fa1_s2_r[20] ,
         \mul_b1/fa1_s2_r[19] , \mul_b1/fa1_s2_r[18] , \mul_b1/fa1_s2_r[17] ,
         \mul_b1/fa1_s2_r[16] , \mul_b1/fa1_s2_r[15] , \mul_b1/fa1_s2_r[14] ,
         \mul_b1/fa1_s2_r[13] , \mul_b1/fa1_c1_r[22] , \mul_b1/fa1_c1_r[21] ,
         \mul_b1/fa1_c1_r[20] , \mul_b1/fa1_c1_r[19] , \mul_b1/fa1_c1_r[18] ,
         \mul_b1/fa1_c1_r[17] , \mul_b1/fa1_c1_r[16] , \mul_b1/fa1_c1_r[15] ,
         \mul_b1/fa1_c1_r[14] , \mul_b1/fa1_c1_r[13] , \mul_b1/fa1_c1_r[12] ,
         \mul_b1/fa1_c1_r[11] , \mul_b1/fa1_c1_r[10] , \mul_b1/fa1_c1_r[9] ,
         \mul_b1/fa1_c1_r[8] , \mul_b1/fa1_s1_r[33] , \mul_b1/fa1_s1_r[32] ,
         \mul_b1/fa1_s1_r[31] , \mul_b1/fa1_s1_r[30] , \mul_b1/fa1_s1_r[29] ,
         \mul_b1/fa1_s1_r[28] , \mul_b1/fa1_s1_r[27] , \mul_b1/fa1_s1_r[26] ,
         \mul_b1/fa1_s1_r[25] , \mul_b1/fa1_s1_r[24] , \mul_b1/fa1_s1_r[23] ,
         \mul_b1/fa1_s1_r[22] , \mul_b1/fa1_s1_r[21] , \mul_b1/fa1_s1_r[20] ,
         \mul_b1/fa1_s1_r[19] , \mul_b1/fa1_s1_r[18] , \mul_b1/fa1_s1_r[17] ,
         \mul_b1/fa1_s1_r[16] , \mul_b1/fa1_s1_r[15] , \mul_b1/fa1_s1_r[14] ,
         \mul_b1/fa1_s1_r[13] , \mul_b1/fa1_s1_r[12] , \mul_b1/fa1_s1_r[11] ,
         \mul_b1/fa1_s1_r[10] , \mul_b1/fa1_s1_r[9] , \mul_b1/fa1_s1_r[8] ,
         \mul_b1/fa1_s1_r[7] , \mul_b1/fa1_s1_r[6] , \mul_b1/fa1_s0_r[33] ,
         \mul_b1/fa1_s0_r[32] , \mul_b1/fa1_s0_r[31] , \mul_b1/fa1_s0_r[30] ,
         \mul_b1/fa1_s0_r[29] , \mul_b1/fa1_s0_r[28] , \mul_b1/fa1_s0_r[27] ,
         \mul_b1/fa1_s0_r[26] , \mul_b1/fa1_s0_r[25] , \mul_b1/fa1_s0_r[24] ,
         \mul_b1/fa1_s0_r[23] , \mul_b1/fa1_s0_r[22] , \mul_b1/fa1_s0_r[21] ,
         \mul_b1/fa1_s0_r[20] , \mul_b1/fa1_s0_r[19] , \mul_b1/fa1_s0_r[18] ,
         \mul_b1/fa1_s0_r[17] , \mul_b1/fa1_s0_r[16] , \mul_b1/fa1_s0_r[15] ,
         \mul_b1/fa1_s0_r[14] , \mul_b1/fa1_s0_r[13] , \mul_b1/fa1_s0_r[12] ,
         \mul_b1/fa1_s0_r[11] , \mul_b1/fa1_s0_r[10] , \mul_b1/fa1_s0_r[9] ,
         \mul_b1/fa1_s0_r[8] , \mul_b1/fa1_s0_r[7] , \mul_b1/fa1_s0_r[6] ,
         \mul_b1/fa1_c2[28] , \mul_b1/fa1_c2[27] , \mul_b1/fa1_c2[26] ,
         \mul_b1/fa1_c2[25] , \mul_b1/fa1_c2[24] , \mul_b1/fa1_c2[23] ,
         \mul_b1/fa1_c2[22] , \mul_b1/fa1_c2[21] , \mul_b1/fa1_c2[20] ,
         \mul_b1/fa1_c2[19] , \mul_b1/fa1_c2[18] , \mul_b1/fa1_c2[17] ,
         \mul_b1/fa1_c2[16] , \mul_b1/fa1_c2[15] , \mul_b1/fa1_c2[14] ,
         \mul_b1/fa1_s2[29] , \mul_b1/fa1_s2[28] , \mul_b1/fa1_s2[27] ,
         \mul_b1/fa1_s2[26] , \mul_b1/fa1_s2[25] , \mul_b1/fa1_s2[24] ,
         \mul_b1/fa1_s2[23] , \mul_b1/fa1_s2[22] , \mul_b1/fa1_s2[21] ,
         \mul_b1/fa1_s2[20] , \mul_b1/fa1_s2[19] , \mul_b1/fa1_s2[18] ,
         \mul_b1/fa1_s2[17] , \mul_b1/fa1_s2[16] , \mul_b1/fa1_s2[15] ,
         \mul_b1/fa1_s2[14] , \mul_b1/fa1_c1[22] , \mul_b1/fa1_c1[21] ,
         \mul_b1/fa1_c1[20] , \mul_b1/fa1_c1[19] , \mul_b1/fa1_c1[18] ,
         \mul_b1/fa1_c1[17] , \mul_b1/fa1_c1[16] , \mul_b1/fa1_c1[15] ,
         \mul_b1/fa1_c1[14] , \mul_b1/fa1_c1[13] , \mul_b1/fa1_c1[12] ,
         \mul_b1/fa1_c1[11] , \mul_b1/fa1_c1[10] , \mul_b1/fa1_c1[9] ,
         \mul_b1/fa1_c1[8] , \mul_b1/fa1_s1[27] , \mul_b1/fa1_s1[22] ,
         \mul_b1/fa1_s1[21] , \mul_b1/fa1_s1[20] , \mul_b1/fa1_s1[19] ,
         \mul_b1/fa1_s1[18] , \mul_b1/fa1_s1[17] , \mul_b1/fa1_s1[16] ,
         \mul_b1/fa1_s1[15] , \mul_b1/fa1_s1[14] , \mul_b1/fa1_s1[13] ,
         \mul_b1/fa1_s1[12] , \mul_b1/fa1_s1[11] , \mul_b1/fa1_s1[10] ,
         \mul_b1/fa1_s1[9] , \mul_b1/fa1_s1[8] , \mul_b1/fa1_s1[7] ,
         \mul_b2/result_sat[15] , \mul_b2/result_sat[14] ,
         \mul_b2/result_sat[13] , \mul_b2/result_sat[12] ,
         \mul_b2/result_sat[11] , \mul_b2/result_sat[10] ,
         \mul_b2/result_sat[9] , \mul_b2/result_sat[8] ,
         \mul_b2/result_sat[7] , \mul_b2/result_sat[6] ,
         \mul_b2/result_sat[5] , \mul_b2/result_sat[4] ,
         \mul_b2/result_sat[3] , \mul_b2/result_sat[2] ,
         \mul_b2/result_sat[1] , \mul_b2/result_sat[0] , \mul_b2/fa1_s2_r[33] ,
         \mul_b2/fa1_s2_r[32] , \mul_b2/fa1_s2_r[31] , \mul_b2/fa1_s2_r[30] ,
         \mul_b2/fa1_s2_r[29] , \mul_b2/fa1_s2_r[28] , \mul_b2/fa1_s2_r[27] ,
         \mul_b2/fa1_s2_r[26] , \mul_b2/fa1_s2_r[25] , \mul_b2/fa1_s2_r[24] ,
         \mul_b2/fa1_s2_r[23] , \mul_b2/fa1_s2_r[22] , \mul_b2/fa1_s2_r[21] ,
         \mul_b2/fa1_s2_r[20] , \mul_b2/fa1_s2_r[19] , \mul_b2/fa1_s2_r[18] ,
         \mul_b2/fa1_s2_r[17] , \mul_b2/fa1_s2_r[16] , \mul_b2/fa1_s2_r[15] ,
         \mul_b2/fa1_s2_r[14] , \mul_b2/fa1_s2_r[13] , \mul_b2/fa1_s2_r[12] ,
         \mul_b2/fa1_s1_r[33] , \mul_b2/fa1_s1_r[32] , \mul_b2/fa1_s1_r[31] ,
         \mul_b2/fa1_s1_r[30] , \mul_b2/fa1_s1_r[29] , \mul_b2/fa1_s1_r[28] ,
         \mul_b2/fa1_s1_r[27] , \mul_b2/fa1_s1_r[26] , \mul_b2/fa1_s1_r[25] ,
         \mul_b2/fa1_s1_r[24] , \mul_b2/fa1_s1_r[23] , \mul_b2/fa1_s1_r[22] ,
         \mul_b2/fa1_s1_r[21] , \mul_b2/fa1_s1_r[20] , \mul_b2/fa1_s1_r[19] ,
         \mul_b2/fa1_s1_r[18] , \mul_b2/fa1_s1_r[17] , \mul_b2/fa1_s1_r[16] ,
         \mul_b2/fa1_s1_r[15] , \mul_b2/fa1_s1_r[14] , \mul_b2/fa1_s1_r[13] ,
         \mul_b2/fa1_s1_r[12] , \mul_b2/fa1_s1_r[11] , \mul_b2/fa1_s1_r[10] ,
         \mul_b2/fa1_s1_r[9] , \mul_b2/fa1_s1_r[8] , \mul_b2/fa1_s1_r[7] ,
         \mul_b2/fa1_s1_r[6] , \mul_b2/fa1_c0_r[32] , \mul_b2/fa1_c0_r[31] ,
         \mul_b2/fa1_c0_r[30] , \mul_b2/fa1_c0_r[29] , \mul_b2/fa1_c0_r[28] ,
         \mul_b2/fa1_c0_r[27] , \mul_b2/fa1_c0_r[26] , \mul_b2/fa1_c0_r[25] ,
         \mul_b2/fa1_c0_r[24] , \mul_b2/fa1_c0_r[23] , \mul_b2/fa1_c0_r[22] ,
         \mul_b2/fa1_c0_r[21] , \mul_b2/fa1_c0_r[20] , \mul_b2/fa1_c0_r[19] ,
         \mul_b2/fa1_c0_r[18] , \mul_b2/fa1_c0_r[17] , \mul_b2/fa1_c0_r[16] ,
         \mul_b2/fa1_c0_r[15] , \mul_b2/fa1_c0_r[14] , \mul_b2/fa1_c0_r[13] ,
         \mul_b2/fa1_c0_r[12] , \mul_b2/fa1_c0_r[11] , \mul_b2/fa1_c0_r[10] ,
         \mul_b2/fa1_c0_r[9] , \mul_b2/fa1_c0_r[8] , \mul_b2/fa1_c0_r[7] ,
         \mul_b2/fa1_c0_r[6] , \mul_b2/fa1_c0_r[5] , \mul_b2/fa1_c0_r[4] ,
         \mul_b2/fa1_s0_r[18] , \mul_b2/fa1_s0_r[17] , \mul_b2/fa1_s0_r[16] ,
         \mul_b2/fa1_s0_r[15] , \mul_b2/fa1_s0_r[14] , \mul_b2/fa1_s0_r[13] ,
         \mul_b2/fa1_s0_r[12] , \mul_b2/fa1_s0_r[11] , \mul_b2/fa1_s0_r[10] ,
         \mul_b2/fa1_s0_r[9] , \mul_b2/fa1_s0_r[8] , \mul_b2/fa1_s0_r[7] ,
         \mul_b2/fa1_s0_r[6] , \mul_b2/fa1_s0_r[5] , \mul_b2/fa1_s1[7] ,
         \mul_b2/fa1_c0[18] , \mul_b2/fa1_c0[17] , \mul_b2/fa1_c0[16] ,
         \mul_b2/fa1_c0[15] , \mul_b2/fa1_c0[14] , \mul_b2/fa1_c0[13] ,
         \mul_b2/fa1_c0[12] , \mul_b2/fa1_c0[11] , \mul_b2/fa1_c0[10] ,
         \mul_b2/fa1_c0[9] , \mul_b2/fa1_c0[8] , \mul_b2/fa1_c0[7] ,
         \mul_b2/fa1_c0[6] , \mul_b2/fa1_c0[5] , \mul_b2/fa1_c0[4] ,
         \mul_b2/fa1_s0[18] , \mul_b2/fa1_s0[17] , \mul_b2/fa1_s0[16] ,
         \mul_b2/fa1_s0[15] , \mul_b2/fa1_s0[14] , \mul_b2/fa1_s0[13] ,
         \mul_b2/fa1_s0[12] , \mul_b2/fa1_s0[11] , \mul_b2/fa1_s0[10] ,
         \mul_b2/fa1_s0[9] , \mul_b2/fa1_s0[8] , \mul_b2/fa1_s0[7] ,
         \mul_b2/fa1_s0[6] , \mul_b2/fa1_s0[5] , \mul_a1/result_sat[15] ,
         \mul_a1/result_sat[14] , \mul_a1/result_sat[13] ,
         \mul_a1/result_sat[12] , \mul_a1/result_sat[11] ,
         \mul_a1/result_sat[10] , \mul_a1/result_sat[9] ,
         \mul_a1/result_sat[8] , \mul_a1/result_sat[7] ,
         \mul_a1/result_sat[6] , \mul_a1/result_sat[5] ,
         \mul_a1/result_sat[4] , \mul_a1/result_sat[3] ,
         \mul_a1/result_sat[2] , \mul_a1/result_sat[1] ,
         \mul_a1/result_sat[0] , \mul_a1/fa1_s2_r[33] , \mul_a1/fa1_s2_r[32] ,
         \mul_a1/fa1_s2_r[31] , \mul_a1/fa1_s2_r[30] , \mul_a1/fa1_s2_r[29] ,
         \mul_a1/fa1_s2_r[28] , \mul_a1/fa1_s2_r[27] , \mul_a1/fa1_s2_r[26] ,
         \mul_a1/fa1_s2_r[25] , \mul_a1/fa1_s2_r[24] , \mul_a1/fa1_s2_r[23] ,
         \mul_a1/fa1_s2_r[22] , \mul_a1/fa1_s2_r[21] , \mul_a1/fa1_s2_r[20] ,
         \mul_a1/fa1_s2_r[19] , \mul_a1/fa1_s2_r[18] , \mul_a1/fa1_s2_r[17] ,
         \mul_a1/fa1_s2_r[16] , \mul_a1/fa1_s2_r[15] , \mul_a1/fa1_s2_r[14] ,
         \mul_a1/fa1_s2_r[13] , \mul_a1/fa1_s2_r[12] , \mul_a1/fa1_c1_r[25] ,
         \mul_a1/fa1_c1_r[24] , \mul_a1/fa1_c1_r[23] , \mul_a1/fa1_c1_r[22] ,
         \mul_a1/fa1_c1_r[21] , \mul_a1/fa1_c1_r[20] , \mul_a1/fa1_c1_r[19] ,
         \mul_a1/fa1_c1_r[18] , \mul_a1/fa1_c1_r[17] , \mul_a1/fa1_c1_r[16] ,
         \mul_a1/fa1_c1_r[15] , \mul_a1/fa1_c1_r[14] , \mul_a1/fa1_c1_r[13] ,
         \mul_a1/fa1_c1_r[12] , \mul_a1/fa1_c1_r[11] , \mul_a1/fa1_s1_r[33] ,
         \mul_a1/fa1_s1_r[32] , \mul_a1/fa1_s1_r[31] , \mul_a1/fa1_s1_r[30] ,
         \mul_a1/fa1_s1_r[29] , \mul_a1/fa1_s1_r[28] , \mul_a1/fa1_s1_r[27] ,
         \mul_a1/fa1_s1_r[26] , \mul_a1/fa1_s1_r[25] , \mul_a1/fa1_s1_r[24] ,
         \mul_a1/fa1_s1_r[23] , \mul_a1/fa1_s1_r[22] , \mul_a1/fa1_s1_r[21] ,
         \mul_a1/fa1_s1_r[20] , \mul_a1/fa1_s1_r[19] , \mul_a1/fa1_s1_r[18] ,
         \mul_a1/fa1_s1_r[17] , \mul_a1/fa1_s1_r[16] , \mul_a1/fa1_s1_r[15] ,
         \mul_a1/fa1_s1_r[14] , \mul_a1/fa1_s1_r[13] , \mul_a1/fa1_s1_r[12] ,
         \mul_a1/fa1_s1_r[11] , \mul_a1/fa1_s1_r[10] , \mul_a1/fa1_s1_r[9] ,
         \mul_a1/fa1_c0_r[17] , \mul_a1/fa1_c0_r[16] , \mul_a1/fa1_c0_r[15] ,
         \mul_a1/fa1_c0_r[14] , \mul_a1/fa1_c0_r[13] , \mul_a1/fa1_c0_r[12] ,
         \mul_a1/fa1_c0_r[11] , \mul_a1/fa1_c0_r[10] , \mul_a1/fa1_c0_r[9] ,
         \mul_a1/fa1_c0_r[8] , \mul_a1/fa1_c0_r[7] , \mul_a1/fa1_c0_r[6] ,
         \mul_a1/fa1_c0_r[5] , \mul_a1/fa1_c0_r[4] , \mul_a1/fa1_c0_r[3] ,
         \mul_a1/fa1_s0_r[33] , \mul_a1/fa1_s0_r[32] , \mul_a1/fa1_s0_r[31] ,
         \mul_a1/fa1_s0_r[30] , \mul_a1/fa1_s0_r[29] , \mul_a1/fa1_s0_r[28] ,
         \mul_a1/fa1_s0_r[27] , \mul_a1/fa1_s0_r[26] , \mul_a1/fa1_s0_r[25] ,
         \mul_a1/fa1_s0_r[24] , \mul_a1/fa1_s0_r[23] , \mul_a1/fa1_s0_r[22] ,
         \mul_a1/fa1_s0_r[21] , \mul_a1/fa1_s0_r[20] , \mul_a1/fa1_s0_r[19] ,
         \mul_a1/fa1_s0_r[18] , \mul_a1/fa1_s0_r[17] , \mul_a1/fa1_s0_r[16] ,
         \mul_a1/fa1_s0_r[15] , \mul_a1/fa1_s0_r[14] , \mul_a1/fa1_s0_r[13] ,
         \mul_a1/fa1_s0_r[12] , \mul_a1/fa1_s0_r[11] , \mul_a1/fa1_s0_r[10] ,
         \mul_a1/fa1_s0_r[9] , \mul_a1/fa1_s0_r[8] , \mul_a1/fa1_s0_r[7] ,
         \mul_a1/fa1_s0_r[6] , \mul_a1/fa1_s0_r[5] , \mul_a1/fa1_s0_r[4] ,
         \mul_a1/fa1_c1[25] , \mul_a1/fa1_c1[24] , \mul_a1/fa1_c1[23] ,
         \mul_a1/fa1_c1[22] , \mul_a1/fa1_c1[21] , \mul_a1/fa1_c1[20] ,
         \mul_a1/fa1_c1[19] , \mul_a1/fa1_c1[18] , \mul_a1/fa1_c1[17] ,
         \mul_a1/fa1_c1[16] , \mul_a1/fa1_c1[15] , \mul_a1/fa1_c1[14] ,
         \mul_a1/fa1_c1[13] , \mul_a1/fa1_c1[12] , \mul_a1/fa1_c1[11] ,
         \mul_a1/fa1_s1[29] , \mul_a1/fa1_s1[25] , \mul_a1/fa1_s1[24] ,
         \mul_a1/fa1_s1[23] , \mul_a1/fa1_s1[22] , \mul_a1/fa1_s1[21] ,
         \mul_a1/fa1_s1[20] , \mul_a1/fa1_s1[19] , \mul_a1/fa1_s1[18] ,
         \mul_a1/fa1_s1[17] , \mul_a1/fa1_s1[16] , \mul_a1/fa1_s1[15] ,
         \mul_a1/fa1_s1[14] , \mul_a1/fa1_s1[13] , \mul_a1/fa1_s1[12] ,
         \mul_a1/fa1_s1[11] , \mul_a1/fa1_c0[17] , \mul_a1/fa1_c0[16] ,
         \mul_a1/fa1_c0[15] , \mul_a1/fa1_c0[14] , \mul_a1/fa1_c0[13] ,
         \mul_a1/fa1_c0[12] , \mul_a1/fa1_c0[11] , \mul_a1/fa1_c0[10] ,
         \mul_a1/fa1_c0[9] , \mul_a1/fa1_c0[8] , \mul_a1/fa1_c0[7] ,
         \mul_a1/fa1_c0[6] , \mul_a1/fa1_c0[5] , \mul_a1/fa1_c0[4] ,
         \mul_a1/fa1_c0[3] , \mul_a1/fa1_s0[29] , \mul_a1/fa1_s0[17] ,
         \mul_a1/fa1_s0[16] , \mul_a1/fa1_s0[15] , \mul_a1/fa1_s0[14] ,
         \mul_a1/fa1_s0[13] , \mul_a1/fa1_s0[12] , \mul_a1/fa1_s0[11] ,
         \mul_a1/fa1_s0[10] , \mul_a1/fa1_s0[9] , \mul_a1/fa1_s0[8] ,
         \mul_a1/fa1_s0[7] , \mul_a1/fa1_s0[6] , \mul_a1/fa1_s0[5] ,
         \mul_a1/fa1_s0[4] , \mul_a2/result_sat[15] , \mul_a2/result_sat[14] ,
         \mul_a2/result_sat[13] , \mul_a2/result_sat[12] ,
         \mul_a2/result_sat[11] , \mul_a2/result_sat[10] ,
         \mul_a2/result_sat[9] , \mul_a2/result_sat[8] ,
         \mul_a2/result_sat[7] , \mul_a2/result_sat[6] ,
         \mul_a2/result_sat[5] , \mul_a2/result_sat[4] ,
         \mul_a2/result_sat[3] , \mul_a2/result_sat[2] ,
         \mul_a2/result_sat[1] , \mul_a2/result_sat[0] , \mul_a2/fa1_c2_r[28] ,
         \mul_a2/fa1_c2_r[27] , \mul_a2/fa1_c2_r[26] , \mul_a2/fa1_c2_r[25] ,
         \mul_a2/fa1_c2_r[24] , \mul_a2/fa1_c2_r[23] , \mul_a2/fa1_c2_r[22] ,
         \mul_a2/fa1_c2_r[21] , \mul_a2/fa1_c2_r[20] , \mul_a2/fa1_c2_r[19] ,
         \mul_a2/fa1_c2_r[18] , \mul_a2/fa1_c2_r[17] , \mul_a2/fa1_c2_r[16] ,
         \mul_a2/fa1_c2_r[15] , \mul_a2/fa1_c2_r[14] , \mul_a2/fa1_s2_r[33] ,
         \mul_a2/fa1_s2_r[32] , \mul_a2/fa1_s2_r[31] , \mul_a2/fa1_s2_r[30] ,
         \mul_a2/fa1_s2_r[29] , \mul_a2/fa1_s2_r[28] , \mul_a2/fa1_s2_r[27] ,
         \mul_a2/fa1_s2_r[26] , \mul_a2/fa1_s2_r[25] , \mul_a2/fa1_s2_r[24] ,
         \mul_a2/fa1_s2_r[23] , \mul_a2/fa1_s2_r[22] , \mul_a2/fa1_s2_r[21] ,
         \mul_a2/fa1_s2_r[20] , \mul_a2/fa1_s2_r[19] , \mul_a2/fa1_s2_r[18] ,
         \mul_a2/fa1_s2_r[17] , \mul_a2/fa1_s2_r[16] , \mul_a2/fa1_s2_r[15] ,
         \mul_a2/fa1_s2_r[14] , \mul_a2/fa1_s2_r[13] , \mul_a2/fa1_s2_r[12] ,
         \mul_a2/fa1_c1_r[32] , \mul_a2/fa1_c1_r[31] , \mul_a2/fa1_c1_r[30] ,
         \mul_a2/fa1_c1_r[29] , \mul_a2/fa1_c1_r[28] , \mul_a2/fa1_c1_r[27] ,
         \mul_a2/fa1_c1_r[26] , \mul_a2/fa1_c1_r[25] , \mul_a2/fa1_c1_r[24] ,
         \mul_a2/fa1_c1_r[23] , \mul_a2/fa1_c1_r[22] , \mul_a2/fa1_c1_r[21] ,
         \mul_a2/fa1_c1_r[20] , \mul_a2/fa1_c1_r[19] , \mul_a2/fa1_c1_r[18] ,
         \mul_a2/fa1_c1_r[17] , \mul_a2/fa1_c1_r[16] , \mul_a2/fa1_c1_r[15] ,
         \mul_a2/fa1_c1_r[14] , \mul_a2/fa1_c1_r[13] , \mul_a2/fa1_c1_r[12] ,
         \mul_a2/fa1_c1_r[11] , \mul_a2/fa1_c1_r[10] , \mul_a2/fa1_c1_r[9] ,
         \mul_a2/fa1_c1_r[8] , \mul_a2/fa1_s1_r[23] , \mul_a2/fa1_s1_r[22] ,
         \mul_a2/fa1_s1_r[21] , \mul_a2/fa1_s1_r[20] , \mul_a2/fa1_s1_r[19] ,
         \mul_a2/fa1_s1_r[18] , \mul_a2/fa1_s1_r[17] , \mul_a2/fa1_s1_r[16] ,
         \mul_a2/fa1_s1_r[15] , \mul_a2/fa1_s1_r[14] , \mul_a2/fa1_s1_r[13] ,
         \mul_a2/fa1_s1_r[12] , \mul_a2/fa1_s1_r[11] , \mul_a2/fa1_s1_r[10] ,
         \mul_a2/fa1_s1_r[9] , \mul_a2/fa1_s1_r[8] , \mul_a2/fa1_s1_r[7] ,
         \mul_a2/fa1_s0_r[33] , \mul_a2/fa1_s0_r[32] , \mul_a2/fa1_s0_r[31] ,
         \mul_a2/fa1_s0_r[30] , \mul_a2/fa1_s0_r[29] , \mul_a2/fa1_s0_r[28] ,
         \mul_a2/fa1_s0_r[27] , \mul_a2/fa1_s0_r[26] , \mul_a2/fa1_s0_r[25] ,
         \mul_a2/fa1_s0_r[24] , \mul_a2/fa1_s0_r[23] , \mul_a2/fa1_s0_r[22] ,
         \mul_a2/fa1_s0_r[21] , \mul_a2/fa1_s0_r[20] , \mul_a2/fa1_s0_r[19] ,
         \mul_a2/fa1_s0_r[18] , \mul_a2/fa1_s0_r[17] , \mul_a2/fa1_s0_r[16] ,
         \mul_a2/fa1_s0_r[15] , \mul_a2/fa1_s0_r[14] , \mul_a2/fa1_s0_r[13] ,
         \mul_a2/fa1_s0_r[12] , \mul_a2/fa1_s0_r[11] , \mul_a2/fa1_s0_r[10] ,
         \mul_a2/fa1_s0_r[9] , \mul_a2/fa1_s0_r[8] , \mul_a2/fa1_s0_r[7] ,
         \mul_a2/fa1_c2[28] , \mul_a2/fa1_c2[27] , \mul_a2/fa1_c2[26] ,
         \mul_a2/fa1_c2[25] , \mul_a2/fa1_c2[24] , \mul_a2/fa1_c2[23] ,
         \mul_a2/fa1_c2[22] , \mul_a2/fa1_c2[21] , \mul_a2/fa1_c2[20] ,
         \mul_a2/fa1_c2[19] , \mul_a2/fa1_c2[18] , \mul_a2/fa1_c2[17] ,
         \mul_a2/fa1_c2[16] , \mul_a2/fa1_c2[15] , \mul_a2/fa1_c2[14] ,
         \mul_a2/fa1_s2[29] , \mul_a2/fa1_s2[28] , \mul_a2/fa1_s2[27] ,
         \mul_a2/fa1_s2[26] , \mul_a2/fa1_s2[25] , \mul_a2/fa1_s2[24] ,
         \mul_a2/fa1_s2[23] , \mul_a2/fa1_s2[22] , \mul_a2/fa1_s2[21] ,
         \mul_a2/fa1_s2[20] , \mul_a2/fa1_s2[19] , \mul_a2/fa1_s2[18] ,
         \mul_a2/fa1_s2[17] , \mul_a2/fa1_s2[16] , \mul_a2/fa1_s2[15] ,
         \mul_a2/fa1_s2[14] , \mul_a2/fa1_c1[24] , \mul_a2/fa1_c1[22] ,
         \mul_a2/fa1_c1[21] , \mul_a2/fa1_c1[20] , \mul_a2/fa1_c1[19] ,
         \mul_a2/fa1_c1[18] , \mul_a2/fa1_c1[17] , \mul_a2/fa1_c1[16] ,
         \mul_a2/fa1_c1[15] , \mul_a2/fa1_c1[14] , \mul_a2/fa1_c1[13] ,
         \mul_a2/fa1_c1[12] , \mul_a2/fa1_c1[11] , \mul_a2/fa1_c1[10] ,
         \mul_a2/fa1_c1[9] , \mul_a2/fa1_c1[8] , \mul_a2/fa1_s1[23] ,
         \mul_a2/fa1_s1[22] , \mul_a2/fa1_s1[21] , \mul_a2/fa1_s1[20] ,
         \mul_a2/fa1_s1[19] , \mul_a2/fa1_s1[18] , \mul_a2/fa1_s1[17] ,
         \mul_a2/fa1_s1[16] , \mul_a2/fa1_s1[15] , \mul_a2/fa1_s1[14] ,
         \mul_a2/fa1_s1[13] , \mul_a2/fa1_s1[12] , \mul_a2/fa1_s1[11] ,
         \mul_a2/fa1_s1[10] , \mul_a2/fa1_s1[9] , \mul_a2/fa1_s1[8] ,
         \C64/DATA4_13 , \C55/DATA4_13 , \C55/DATA4_14 , \C55/DATA4_15 ,
         \C55/DATA4_16 , \C55/DATA4_17 , \C55/DATA4_18 , \C55/DATA4_19 ,
         \C55/DATA4_20 , \C55/DATA4_21 , \C55/DATA4_22 , \C55/DATA4_23 ,
         \C55/DATA4_24 , \C55/DATA4_25 , \C55/DATA4_26 , \C55/DATA4_27 ,
         \C55/DATA4_28 , \C53/DATA4_10 , \C43/DATA4_8 , \C43/DATA4_9 ,
         \C43/DATA4_10 , \C43/DATA4_11 , \C43/DATA4_12 , \C43/DATA4_13 ,
         \C43/DATA4_14 , \C43/DATA4_15 , \C43/DATA4_16 , \C43/DATA4_17 ,
         \C43/DATA4_18 , \C43/DATA4_19 , \C43/DATA4_20 , \C43/DATA4_21 ,
         \C43/DATA4_22 , \C33/DATA4_6 , \C33/DATA4_7 , \C33/DATA4_8 ,
         \C33/DATA4_9 , \C33/DATA4_10 , \C33/DATA4_11 , \C33/DATA4_12 ,
         \C33/DATA4_13 , \C33/DATA4_14 , \C33/DATA4_15 , \C33/DATA4_16 ,
         \C33/DATA4_17 , \C33/DATA4_18 , \C33/DATA4_19 , \C33/DATA4_20 , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888;
  wire   [15:0] x_z1;
  wire   [15:0] x_z2;
  wire   [15:0] y_z1;
  wire   [15:0] y_z2;
  wire   [15:0] x_reg2;
  wire   [15:0] p_b0;
  wire   [15:0] p_b1;
  wire   [15:0] p_b2;
  wire   [15:0] p_a1;
  wire   [15:0] p_a2;

  HS65_GS_DFPRQX4 valid_T1_reg ( .D(n1792), .CP(clk), .RN(rst_n), .Q(valid_T1)
         );
  HS65_GS_DFPRQX4 valid_T2_reg ( .D(valid_T1), .CP(clk), .RN(rst_n), .Q(
        valid_T2) );
  HS65_GS_DFPRQX4 valid_T3_reg ( .D(valid_T2), .CP(clk), .RN(rst_n), .Q(
        valid_T3) );
  HS65_GS_DFPRQX4 valid_out_reg ( .D(valid_T3), .CP(clk), .RN(rst_n), .Q(
        valid_out) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[0]  ( .D(\mul_b0/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[0]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[1]  ( .D(\mul_b0/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[1]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[2]  ( .D(\mul_b0/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[2]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[3]  ( .D(\mul_b0/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[3]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[4]  ( .D(\mul_b0/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[4]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[5]  ( .D(\mul_b0/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[5]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[6]  ( .D(\mul_b0/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[6]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[7]  ( .D(\mul_b0/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[7]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[8]  ( .D(\mul_b0/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[8]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[9]  ( .D(\mul_b0/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[9]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[10]  ( .D(\mul_b0/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[10]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[11]  ( .D(\mul_b0/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[11]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[12]  ( .D(\mul_b0/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[12]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[13]  ( .D(\mul_b0/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[13]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[14]  ( .D(\mul_b0/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[14]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[15]  ( .D(\mul_b0/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[15]) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[12]  ( .D(x_z1[0]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[13]  ( .D(x_z1[1]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[14]  ( .D(x_z1[2]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[15]  ( .D(x_z1[3]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[16]  ( .D(x_z1[4]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[17]  ( .D(x_z1[5]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[18]  ( .D(x_z1[6]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[19]  ( .D(x_z1[7]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[20]  ( .D(x_z1[8]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[21]  ( .D(x_z1[9]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[22]  ( .D(x_z1[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[23]  ( .D(x_z1[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[24]  ( .D(x_z1[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[25]  ( .D(x_z1[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[26]  ( .D(x_z1[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[27]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[28]  ( .D(n1791), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[29]  ( .D(n1791), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[30]  ( .D(n1791), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[31]  ( .D(n1791), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[32]  ( .D(n1791), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[33]  ( .D(n1791), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[8]  ( .D(x_z1[0]), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[9]  ( .D(x_z1[1]), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[10]  ( .D(x_z1[2]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[11]  ( .D(x_z1[3]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[12]  ( .D(x_z1[4]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[13]  ( .D(x_z1[5]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[14]  ( .D(x_z1[6]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[15]  ( .D(x_z1[7]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[16]  ( .D(x_z1[8]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[17]  ( .D(x_z1[9]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[18]  ( .D(x_z1[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[19]  ( .D(x_z1[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[20]  ( .D(x_z1[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[21]  ( .D(x_z1[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[22]  ( .D(x_z1[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[23]  ( .D(n1791), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[24]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[25]  ( .D(n1791), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[26]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[27]  ( .D(n1791), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[28]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[29]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[30]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[31]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[32]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[33]  ( .D(n1791), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[5]  ( .D(\mul_b0/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[6]  ( .D(\mul_b0/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[7]  ( .D(\mul_b0/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[8]  ( .D(\mul_b0/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[9]  ( .D(\mul_b0/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[10]  ( .D(\mul_b0/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[11]  ( .D(\mul_b0/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[12]  ( .D(\mul_b0/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[13]  ( .D(\mul_b0/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[14]  ( .D(\mul_b0/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[15]  ( .D(\mul_b0/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[16]  ( .D(\mul_b0/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[17]  ( .D(\mul_b0/fa1_c0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[18]  ( .D(\mul_b0/fa1_c0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[19]  ( .D(\mul_b0/fa1_c0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[20]  ( .D(\mul_b0/fa1_c0[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[6]  ( .D(\mul_b0/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[7]  ( .D(\mul_b0/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[8]  ( .D(\mul_b0/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[9]  ( .D(\mul_b0/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[10]  ( .D(\mul_b0/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[11]  ( .D(\mul_b0/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[12]  ( .D(\mul_b0/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[13]  ( .D(\mul_b0/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[14]  ( .D(\mul_b0/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[15]  ( .D(\mul_b0/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[16]  ( .D(\mul_b0/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[17]  ( .D(\mul_b0/fa1_s0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[18]  ( .D(\mul_b0/fa1_s0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[19]  ( .D(\mul_b0/fa1_s0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[20]  ( .D(\mul_b0/fa1_s0[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[21]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[22]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[23]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[24]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[25]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[26]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[27]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[28]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[29]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[30]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[31]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[32]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[33]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[0]  ( .D(\mul_b1/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[0]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[1]  ( .D(\mul_b1/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[1]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[2]  ( .D(\mul_b1/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[2]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[3]  ( .D(\mul_b1/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[3]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[4]  ( .D(\mul_b1/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[4]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[5]  ( .D(\mul_b1/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[5]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[6]  ( .D(\mul_b1/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[6]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[7]  ( .D(\mul_b1/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[7]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[8]  ( .D(\mul_b1/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[8]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[9]  ( .D(\mul_b1/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[9]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[10]  ( .D(\mul_b1/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[10]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[11]  ( .D(\mul_b1/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[11]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[12]  ( .D(\mul_b1/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[12]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[13]  ( .D(\mul_b1/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[13]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[14]  ( .D(\mul_b1/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[14]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[15]  ( .D(\mul_b1/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[15]) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[13]  ( .D(x_z2[0]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[14]  ( .D(\mul_b1/fa1_s2[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[15]  ( .D(\mul_b1/fa1_s2[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[16]  ( .D(\mul_b1/fa1_s2[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[17]  ( .D(\mul_b1/fa1_s2[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[18]  ( .D(\mul_b1/fa1_s2[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[19]  ( .D(\mul_b1/fa1_s2[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[20]  ( .D(\mul_b1/fa1_s2[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[21]  ( .D(\mul_b1/fa1_s2[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[22]  ( .D(\mul_b1/fa1_s2[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[23]  ( .D(\mul_b1/fa1_s2[23] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[24]  ( .D(\mul_b1/fa1_s2[24] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[25]  ( .D(\mul_b1/fa1_s2[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[26]  ( .D(\mul_b1/fa1_s2[26] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[27]  ( .D(\mul_b1/fa1_s2[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[28]  ( .D(\mul_b1/fa1_s2[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[29]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[30]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[31]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[32]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[33]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[8]  ( .D(\mul_b1/fa1_c1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[9]  ( .D(\mul_b1/fa1_c1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[10]  ( .D(\mul_b1/fa1_c1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[11]  ( .D(\mul_b1/fa1_c1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[12]  ( .D(\mul_b1/fa1_c1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[13]  ( .D(\mul_b1/fa1_c1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[14]  ( .D(\mul_b1/fa1_c1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[15]  ( .D(\mul_b1/fa1_c1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[16]  ( .D(\mul_b1/fa1_c1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[17]  ( .D(\mul_b1/fa1_c1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[18]  ( .D(\mul_b1/fa1_c1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[19]  ( .D(\mul_b1/fa1_c1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[20]  ( .D(\mul_b1/fa1_c1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[21]  ( .D(\mul_b1/fa1_c1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[22]  ( .D(\mul_b1/fa1_c1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[6]  ( .D(x_z2[0]), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s1_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[7]  ( .D(\mul_b1/fa1_s1[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s1_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[8]  ( .D(\mul_b1/fa1_s1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[9]  ( .D(\mul_b1/fa1_s1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[10]  ( .D(\mul_b1/fa1_s1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[11]  ( .D(\mul_b1/fa1_s1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[12]  ( .D(\mul_b1/fa1_s1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[13]  ( .D(\mul_b1/fa1_s1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[14]  ( .D(\mul_b1/fa1_s1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[15]  ( .D(\mul_b1/fa1_s1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[16]  ( .D(\mul_b1/fa1_s1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[17]  ( .D(\mul_b1/fa1_s1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[18]  ( .D(\mul_b1/fa1_s1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[19]  ( .D(\mul_b1/fa1_s1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[20]  ( .D(\mul_b1/fa1_s1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[21]  ( .D(\mul_b1/fa1_s1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[22]  ( .D(\mul_b1/fa1_s1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[23]  ( .D(\mul_b1/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[24]  ( .D(\mul_b1/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[25]  ( .D(\mul_b1/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[26]  ( .D(\mul_b1/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[27]  ( .D(\mul_b1/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[28]  ( .D(\mul_b1/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[29]  ( .D(\mul_b1/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[30]  ( .D(\mul_b1/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[31]  ( .D(\mul_b1/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[32]  ( .D(\mul_b1/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[33]  ( .D(\mul_b1/fa1_s1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[6]  ( .D(\C33/DATA4_6 ), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[7]  ( .D(\C33/DATA4_7 ), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[8]  ( .D(\C33/DATA4_8 ), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[9]  ( .D(\C33/DATA4_9 ), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[10]  ( .D(\C33/DATA4_10 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[11]  ( .D(\C33/DATA4_11 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[12]  ( .D(\C33/DATA4_12 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[13]  ( .D(\C33/DATA4_13 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[14]  ( .D(\C33/DATA4_14 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[15]  ( .D(\C33/DATA4_15 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[16]  ( .D(\C33/DATA4_16 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[17]  ( .D(\C33/DATA4_17 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[18]  ( .D(\C33/DATA4_18 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[19]  ( .D(\C33/DATA4_19 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[20]  ( .D(\C33/DATA4_20 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[21]  ( .D(n1787), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[22]  ( .D(n1787), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[23]  ( .D(n1787), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[24]  ( .D(n1787), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[25]  ( .D(n1787), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[26]  ( .D(n1787), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[27]  ( .D(n1787), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[28]  ( .D(n1787), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[29]  ( .D(n1787), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[30]  ( .D(n1787), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[31]  ( .D(n1787), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[32]  ( .D(n1787), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[33]  ( .D(n1787), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[14]  ( .D(\mul_b1/fa1_c2[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[15]  ( .D(\mul_b1/fa1_c2[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[16]  ( .D(\mul_b1/fa1_c2[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[17]  ( .D(\mul_b1/fa1_c2[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[18]  ( .D(\mul_b1/fa1_c2[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[19]  ( .D(\mul_b1/fa1_c2[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[20]  ( .D(\mul_b1/fa1_c2[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[21]  ( .D(\mul_b1/fa1_c2[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[22]  ( .D(\mul_b1/fa1_c2[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[23]  ( .D(\mul_b1/fa1_c2[23] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[24]  ( .D(\mul_b1/fa1_c2[24] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[25]  ( .D(\mul_b1/fa1_c2[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[26]  ( .D(\mul_b1/fa1_c2[26] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[27]  ( .D(\mul_b1/fa1_c2[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[28]  ( .D(\mul_b1/fa1_c2[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[0]  ( .D(\mul_b2/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[0]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[1]  ( .D(\mul_b2/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[1]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[2]  ( .D(\mul_b2/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[2]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[3]  ( .D(\mul_b2/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[3]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[4]  ( .D(\mul_b2/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[4]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[5]  ( .D(\mul_b2/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[5]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[6]  ( .D(\mul_b2/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[6]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[7]  ( .D(\mul_b2/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[7]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[8]  ( .D(\mul_b2/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[8]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[9]  ( .D(\mul_b2/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[9]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[10]  ( .D(\mul_b2/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[10]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[11]  ( .D(\mul_b2/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[11]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[12]  ( .D(\mul_b2/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[12]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[13]  ( .D(\mul_b2/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[13]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[14]  ( .D(\mul_b2/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[14]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[15]  ( .D(\mul_b2/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[15]) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[12]  ( .D(x_reg2[0]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[13]  ( .D(x_reg2[1]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[14]  ( .D(x_reg2[2]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[15]  ( .D(x_reg2[3]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[16]  ( .D(x_reg2[4]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[17]  ( .D(x_reg2[5]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[18]  ( .D(x_reg2[6]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[19]  ( .D(x_reg2[7]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[20]  ( .D(x_reg2[8]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[21]  ( .D(x_reg2[9]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[22]  ( .D(x_reg2[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[23]  ( .D(x_reg2[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[24]  ( .D(x_reg2[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[25]  ( .D(x_reg2[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[26]  ( .D(x_reg2[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[27]  ( .D(n1789), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[28]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[29]  ( .D(n1789), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[30]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[31]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[32]  ( .D(n1789), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[33]  ( .D(n1789), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[6]  ( .D(x_reg2[0]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[7]  ( .D(\mul_b2/fa1_s1[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[8]  ( .D(\C43/DATA4_8 ), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[9]  ( .D(\C43/DATA4_9 ), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[10]  ( .D(\C43/DATA4_10 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[11]  ( .D(\C43/DATA4_11 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[12]  ( .D(\C43/DATA4_12 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[13]  ( .D(\C43/DATA4_13 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[14]  ( .D(\C43/DATA4_14 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[15]  ( .D(\C43/DATA4_15 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[16]  ( .D(\C43/DATA4_16 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[17]  ( .D(\C43/DATA4_17 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[18]  ( .D(\C43/DATA4_18 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[19]  ( .D(\C43/DATA4_19 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[20]  ( .D(\C43/DATA4_20 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[21]  ( .D(\C43/DATA4_21 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[22]  ( .D(\C43/DATA4_22 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[23]  ( .D(n1786), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[24]  ( .D(n1786), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[25]  ( .D(n1786), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[26]  ( .D(n1786), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[27]  ( .D(n1786), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[28]  ( .D(n1786), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[29]  ( .D(n1786), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[30]  ( .D(n1786), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[31]  ( .D(n1786), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[32]  ( .D(n1786), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[33]  ( .D(n1786), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[4]  ( .D(\mul_b2/fa1_c0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[5]  ( .D(\mul_b2/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[6]  ( .D(\mul_b2/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[7]  ( .D(\mul_b2/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[8]  ( .D(\mul_b2/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[9]  ( .D(\mul_b2/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[10]  ( .D(\mul_b2/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[11]  ( .D(\mul_b2/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[12]  ( .D(\mul_b2/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[13]  ( .D(\mul_b2/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[14]  ( .D(\mul_b2/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[15]  ( .D(\mul_b2/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[16]  ( .D(\mul_b2/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[17]  ( .D(\mul_b2/fa1_c0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[18]  ( .D(\mul_b2/fa1_c0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_c0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[19]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[20]  ( .D(n1789), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[21]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[22]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[23]  ( .D(n1789), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[24]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[25]  ( .D(n1789), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[26]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[27]  ( .D(n1789), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[28]  ( .D(n1789), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[29]  ( .D(n1789), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[30]  ( .D(n1789), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[31]  ( .D(n1789), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_c0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_c0_r_reg[32]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_c0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[5]  ( .D(\mul_b2/fa1_s0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[6]  ( .D(\mul_b2/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[7]  ( .D(\mul_b2/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[8]  ( .D(\mul_b2/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[9]  ( .D(\mul_b2/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[10]  ( .D(\mul_b2/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[11]  ( .D(\mul_b2/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[12]  ( .D(\mul_b2/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[13]  ( .D(\mul_b2/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[14]  ( .D(\mul_b2/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[15]  ( .D(\mul_b2/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[16]  ( .D(\mul_b2/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[17]  ( .D(\mul_b2/fa1_s0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[18]  ( .D(\mul_b2/fa1_s0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b2/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[0]  ( .D(\mul_a1/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[0]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[1]  ( .D(\mul_a1/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[1]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[2]  ( .D(\mul_a1/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[2]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[3]  ( .D(\mul_a1/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[3]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[4]  ( .D(\mul_a1/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[4]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[5]  ( .D(\mul_a1/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[5]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[6]  ( .D(\mul_a1/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[6]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[7]  ( .D(\mul_a1/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[7]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[8]  ( .D(\mul_a1/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[8]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[9]  ( .D(\mul_a1/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[9]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[10]  ( .D(\mul_a1/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[10]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[11]  ( .D(\mul_a1/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[11]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[12]  ( .D(\mul_a1/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[12]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[13]  ( .D(\mul_a1/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[13]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[14]  ( .D(\mul_a1/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[14]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[15]  ( .D(\mul_a1/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[15]) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[12]  ( .D(y_z1[0]), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[13]  ( .D(\C55/DATA4_13 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[14]  ( .D(\C55/DATA4_14 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[15]  ( .D(\C55/DATA4_15 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[16]  ( .D(\C55/DATA4_16 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[17]  ( .D(\C55/DATA4_17 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[18]  ( .D(\C55/DATA4_18 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[19]  ( .D(\C55/DATA4_19 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[20]  ( .D(\C55/DATA4_20 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[21]  ( .D(\C55/DATA4_21 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[22]  ( .D(\C55/DATA4_22 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[23]  ( .D(\C55/DATA4_23 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[24]  ( .D(\C55/DATA4_24 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[25]  ( .D(\C55/DATA4_25 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[26]  ( .D(\C55/DATA4_26 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[27]  ( .D(\C55/DATA4_27 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[28]  ( .D(\C55/DATA4_28 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[29]  ( .D(n1788), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[30]  ( .D(n1788), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[31]  ( .D(n1788), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[32]  ( .D(n1788), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[33]  ( .D(n1788), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[11]  ( .D(\mul_a1/fa1_c1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[12]  ( .D(\mul_a1/fa1_c1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[13]  ( .D(\mul_a1/fa1_c1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[14]  ( .D(\mul_a1/fa1_c1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[15]  ( .D(\mul_a1/fa1_c1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[16]  ( .D(\mul_a1/fa1_c1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[17]  ( .D(\mul_a1/fa1_c1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[18]  ( .D(\mul_a1/fa1_c1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[19]  ( .D(\mul_a1/fa1_c1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[20]  ( .D(\mul_a1/fa1_c1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[21]  ( .D(\mul_a1/fa1_c1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[22]  ( .D(\mul_a1/fa1_c1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[23]  ( .D(\mul_a1/fa1_c1[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[24]  ( .D(\mul_a1/fa1_c1[24] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[25]  ( .D(\mul_a1/fa1_c1[25] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[9]  ( .D(y_z1[0]), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[10]  ( .D(\C53/DATA4_10 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[11]  ( .D(\mul_a1/fa1_s1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[12]  ( .D(\mul_a1/fa1_s1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[13]  ( .D(\mul_a1/fa1_s1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[14]  ( .D(\mul_a1/fa1_s1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[15]  ( .D(\mul_a1/fa1_s1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[16]  ( .D(\mul_a1/fa1_s1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[17]  ( .D(\mul_a1/fa1_s1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[18]  ( .D(\mul_a1/fa1_s1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[19]  ( .D(\mul_a1/fa1_s1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[20]  ( .D(\mul_a1/fa1_s1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[21]  ( .D(\mul_a1/fa1_s1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[22]  ( .D(\mul_a1/fa1_s1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[23]  ( .D(\mul_a1/fa1_s1[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[24]  ( .D(\mul_a1/fa1_s1[24] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[25]  ( .D(\mul_a1/fa1_s1[25] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[26]  ( .D(\mul_a1/fa1_s1[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[27]  ( .D(\mul_a1/fa1_s1[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[28]  ( .D(\mul_a1/fa1_s1[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[29]  ( .D(\mul_a1/fa1_s1[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[30]  ( .D(\mul_a1/fa1_s1[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[31]  ( .D(\mul_a1/fa1_s1[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[32]  ( .D(\mul_a1/fa1_s1[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[33]  ( .D(\mul_a1/fa1_s1[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[3]  ( .D(\mul_a1/fa1_c0[3] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_c0_r[3] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[4]  ( .D(\mul_a1/fa1_c0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_c0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[5]  ( .D(\mul_a1/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[6]  ( .D(\mul_a1/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[7]  ( .D(\mul_a1/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[8]  ( .D(\mul_a1/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[9]  ( .D(\mul_a1/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[10]  ( .D(\mul_a1/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[11]  ( .D(\mul_a1/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[12]  ( .D(\mul_a1/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[13]  ( .D(\mul_a1/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[14]  ( .D(\mul_a1/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[15]  ( .D(\mul_a1/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[16]  ( .D(\mul_a1/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c0_r_reg[17]  ( .D(\mul_a1/fa1_c0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[4]  ( .D(\mul_a1/fa1_s0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[5]  ( .D(\mul_a1/fa1_s0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[6]  ( .D(\mul_a1/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[7]  ( .D(\mul_a1/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[8]  ( .D(\mul_a1/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[9]  ( .D(\mul_a1/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[10]  ( .D(\mul_a1/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[11]  ( .D(\mul_a1/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[12]  ( .D(\mul_a1/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[13]  ( .D(\mul_a1/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[14]  ( .D(\mul_a1/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[15]  ( .D(\mul_a1/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[16]  ( .D(\mul_a1/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[17]  ( .D(\mul_a1/fa1_s0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[18]  ( .D(\mul_a1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[19]  ( .D(\mul_a1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[20]  ( .D(\mul_a1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[21]  ( .D(\mul_a1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[22]  ( .D(\mul_a1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[23]  ( .D(\mul_a1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[24]  ( .D(\mul_a1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[25]  ( .D(\mul_a1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[26]  ( .D(\mul_a1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[27]  ( .D(\mul_a1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[28]  ( .D(\mul_a1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[29]  ( .D(\mul_a1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[30]  ( .D(\mul_a1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[31]  ( .D(\mul_a1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[32]  ( .D(\mul_a1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[33]  ( .D(\mul_a1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[0]  ( .D(\mul_a2/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[0]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[1]  ( .D(\mul_a2/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[1]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[2]  ( .D(\mul_a2/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[2]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[3]  ( .D(\mul_a2/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[3]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[4]  ( .D(\mul_a2/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[4]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[5]  ( .D(\mul_a2/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[5]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[6]  ( .D(\mul_a2/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[6]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[7]  ( .D(\mul_a2/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[7]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[8]  ( .D(\mul_a2/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[8]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[9]  ( .D(\mul_a2/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[9]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[10]  ( .D(\mul_a2/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[10]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[11]  ( .D(\mul_a2/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[11]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[12]  ( .D(\mul_a2/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[12]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[13]  ( .D(\mul_a2/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[13]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[14]  ( .D(\mul_a2/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[14]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[15]  ( .D(\mul_a2/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[15]) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[12]  ( .D(y_z2[0]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[13]  ( .D(\C64/DATA4_13 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[14]  ( .D(\mul_a2/fa1_s2[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[15]  ( .D(\mul_a2/fa1_s2[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[16]  ( .D(\mul_a2/fa1_s2[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[17]  ( .D(\mul_a2/fa1_s2[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[18]  ( .D(\mul_a2/fa1_s2[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[19]  ( .D(\mul_a2/fa1_s2[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[20]  ( .D(\mul_a2/fa1_s2[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[21]  ( .D(\mul_a2/fa1_s2[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[22]  ( .D(\mul_a2/fa1_s2[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[23]  ( .D(\mul_a2/fa1_s2[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[24]  ( .D(\mul_a2/fa1_s2[24] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[25]  ( .D(\mul_a2/fa1_s2[25] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[26]  ( .D(\mul_a2/fa1_s2[26] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[27]  ( .D(\mul_a2/fa1_s2[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[28]  ( .D(\mul_a2/fa1_s2[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[29]  ( .D(\mul_a2/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[30]  ( .D(\mul_a2/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[31]  ( .D(\mul_a2/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[32]  ( .D(\mul_a2/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[33]  ( .D(\mul_a2/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[8]  ( .D(\mul_a2/fa1_c1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[9]  ( .D(\mul_a2/fa1_c1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[10]  ( .D(\mul_a2/fa1_c1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[11]  ( .D(\mul_a2/fa1_c1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[12]  ( .D(\mul_a2/fa1_c1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[13]  ( .D(\mul_a2/fa1_c1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[14]  ( .D(\mul_a2/fa1_c1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[15]  ( .D(\mul_a2/fa1_c1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[16]  ( .D(\mul_a2/fa1_c1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[17]  ( .D(\mul_a2/fa1_c1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[18]  ( .D(\mul_a2/fa1_c1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[19]  ( .D(\mul_a2/fa1_c1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[20]  ( .D(\mul_a2/fa1_c1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[21]  ( .D(\mul_a2/fa1_c1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[22]  ( .D(\mul_a2/fa1_c1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[23]  ( .D(n1785), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[24]  ( .D(\mul_a2/fa1_c1[24] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[25]  ( .D(n1785), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[26]  ( .D(n1785), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[27]  ( .D(n1785), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[28]  ( .D(n1785), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[29]  ( .D(n1785), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[30]  ( .D(n1785), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[31]  ( .D(n1785), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[32]  ( .D(n1785), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[7]  ( .D(y_z2[0]), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s1_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[8]  ( .D(\mul_a2/fa1_s1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[9]  ( .D(\mul_a2/fa1_s1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[10]  ( .D(\mul_a2/fa1_s1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[11]  ( .D(\mul_a2/fa1_s1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[12]  ( .D(\mul_a2/fa1_s1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[13]  ( .D(\mul_a2/fa1_s1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[14]  ( .D(\mul_a2/fa1_s1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[15]  ( .D(\mul_a2/fa1_s1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[16]  ( .D(\mul_a2/fa1_s1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[17]  ( .D(\mul_a2/fa1_s1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[18]  ( .D(\mul_a2/fa1_s1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[19]  ( .D(\mul_a2/fa1_s1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[20]  ( .D(\mul_a2/fa1_s1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[21]  ( .D(\mul_a2/fa1_s1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[22]  ( .D(\mul_a2/fa1_s1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[23]  ( .D(\mul_a2/fa1_s1[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[7]  ( .D(y_z2[7]), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[8]  ( .D(y_z2[8]), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[9]  ( .D(y_z2[9]), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[10]  ( .D(y_z2[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[11]  ( .D(y_z2[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[12]  ( .D(y_z2[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[13]  ( .D(y_z2[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[14]  ( .D(y_z2[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[15]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[16]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[17]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[18]  ( .D(n1790), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[19]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[20]  ( .D(n1790), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[21]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[22]  ( .D(n1790), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[23]  ( .D(n1790), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[24]  ( .D(n1790), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[25]  ( .D(n1790), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[26]  ( .D(n1790), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[27]  ( .D(n1790), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[28]  ( .D(n1790), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[29]  ( .D(n1790), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[30]  ( .D(n1790), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[31]  ( .D(n1790), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[32]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[33]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[14]  ( .D(\mul_a2/fa1_c2[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[15]  ( .D(\mul_a2/fa1_c2[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[16]  ( .D(\mul_a2/fa1_c2[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[17]  ( .D(\mul_a2/fa1_c2[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[18]  ( .D(\mul_a2/fa1_c2[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[19]  ( .D(\mul_a2/fa1_c2[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[20]  ( .D(\mul_a2/fa1_c2[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[21]  ( .D(\mul_a2/fa1_c2[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[22]  ( .D(\mul_a2/fa1_c2[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[23]  ( .D(\mul_a2/fa1_c2[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[24]  ( .D(\mul_a2/fa1_c2[24] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[25]  ( .D(\mul_a2/fa1_c2[25] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[26]  ( .D(\mul_a2/fa1_c2[26] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[27]  ( .D(\mul_a2/fa1_c2[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c2_r_reg[28]  ( .D(\mul_a2/fa1_c2[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c2_r[28] ) );
  HS65_GS_DFPRQX4 \x_z1_reg[15]  ( .D(n1793), .CP(clk), .RN(rst_n), .Q(
        x_z1[15]) );
  HS65_GS_DFPRQX4 \x_z1_reg[14]  ( .D(n1794), .CP(clk), .RN(rst_n), .Q(
        x_z1[14]) );
  HS65_GS_DFPRQX4 \x_z1_reg[13]  ( .D(n1795), .CP(clk), .RN(rst_n), .Q(
        x_z1[13]) );
  HS65_GS_DFPRQX4 \x_z1_reg[12]  ( .D(n1796), .CP(clk), .RN(rst_n), .Q(
        x_z1[12]) );
  HS65_GS_DFPRQX4 \x_z1_reg[11]  ( .D(n1797), .CP(clk), .RN(rst_n), .Q(
        x_z1[11]) );
  HS65_GS_DFPRQX4 \x_z1_reg[10]  ( .D(n1798), .CP(clk), .RN(rst_n), .Q(
        x_z1[10]) );
  HS65_GS_DFPRQX4 \x_z1_reg[9]  ( .D(n1799), .CP(clk), .RN(rst_n), .Q(x_z1[9])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[8]  ( .D(n1800), .CP(clk), .RN(rst_n), .Q(x_z1[8])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[7]  ( .D(n1801), .CP(clk), .RN(rst_n), .Q(x_z1[7])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[6]  ( .D(n1802), .CP(clk), .RN(rst_n), .Q(x_z1[6])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[5]  ( .D(n1803), .CP(clk), .RN(rst_n), .Q(x_z1[5])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[4]  ( .D(n1804), .CP(clk), .RN(rst_n), .Q(x_z1[4])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[3]  ( .D(n1805), .CP(clk), .RN(rst_n), .Q(x_z1[3])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[2]  ( .D(n1806), .CP(clk), .RN(rst_n), .Q(x_z1[2])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[1]  ( .D(n1807), .CP(clk), .RN(rst_n), .Q(x_z1[1])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[0]  ( .D(n1808), .CP(clk), .RN(rst_n), .Q(x_z1[0])
         );
  HS65_GS_DFPRQX4 \x_z2_reg[15]  ( .D(n1809), .CP(clk), .RN(rst_n), .Q(
        x_z2[15]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[15]  ( .D(n1810), .CP(clk), .RN(rst_n), .Q(
        x_reg2[15]) );
  HS65_GS_DFPRQX4 \x_z2_reg[14]  ( .D(n1811), .CP(clk), .RN(rst_n), .Q(
        x_z2[14]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[14]  ( .D(n1812), .CP(clk), .RN(rst_n), .Q(
        x_reg2[14]) );
  HS65_GS_DFPRQX4 \x_z2_reg[13]  ( .D(n1813), .CP(clk), .RN(rst_n), .Q(
        x_z2[13]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[13]  ( .D(n1814), .CP(clk), .RN(rst_n), .Q(
        x_reg2[13]) );
  HS65_GS_DFPRQX4 \x_z2_reg[12]  ( .D(n1815), .CP(clk), .RN(rst_n), .Q(
        x_z2[12]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[12]  ( .D(n1816), .CP(clk), .RN(rst_n), .Q(
        x_reg2[12]) );
  HS65_GS_DFPRQX4 \x_z2_reg[11]  ( .D(n1817), .CP(clk), .RN(rst_n), .Q(
        x_z2[11]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[11]  ( .D(n1818), .CP(clk), .RN(rst_n), .Q(
        x_reg2[11]) );
  HS65_GS_DFPRQX4 \x_z2_reg[10]  ( .D(n1819), .CP(clk), .RN(rst_n), .Q(
        x_z2[10]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[10]  ( .D(n1820), .CP(clk), .RN(rst_n), .Q(
        x_reg2[10]) );
  HS65_GS_DFPRQX4 \x_z2_reg[9]  ( .D(n1821), .CP(clk), .RN(rst_n), .Q(x_z2[9])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[9]  ( .D(n1822), .CP(clk), .RN(rst_n), .Q(
        x_reg2[9]) );
  HS65_GS_DFPRQX4 \x_z2_reg[8]  ( .D(n1823), .CP(clk), .RN(rst_n), .Q(x_z2[8])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[8]  ( .D(n1824), .CP(clk), .RN(rst_n), .Q(
        x_reg2[8]) );
  HS65_GS_DFPRQX4 \x_z2_reg[7]  ( .D(n1825), .CP(clk), .RN(rst_n), .Q(x_z2[7])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[7]  ( .D(n1826), .CP(clk), .RN(rst_n), .Q(
        x_reg2[7]) );
  HS65_GS_DFPRQX4 \x_z2_reg[6]  ( .D(n1827), .CP(clk), .RN(rst_n), .Q(x_z2[6])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[6]  ( .D(n1828), .CP(clk), .RN(rst_n), .Q(
        x_reg2[6]) );
  HS65_GS_DFPRQX4 \x_z2_reg[5]  ( .D(n1829), .CP(clk), .RN(rst_n), .Q(x_z2[5])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[5]  ( .D(n1830), .CP(clk), .RN(rst_n), .Q(
        x_reg2[5]) );
  HS65_GS_DFPRQX4 \x_z2_reg[4]  ( .D(n1831), .CP(clk), .RN(rst_n), .Q(x_z2[4])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[4]  ( .D(n1832), .CP(clk), .RN(rst_n), .Q(
        x_reg2[4]) );
  HS65_GS_DFPRQX4 \x_z2_reg[3]  ( .D(n1833), .CP(clk), .RN(rst_n), .Q(x_z2[3])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[3]  ( .D(n1834), .CP(clk), .RN(rst_n), .Q(
        x_reg2[3]) );
  HS65_GS_DFPRQX4 \x_z2_reg[2]  ( .D(n1835), .CP(clk), .RN(rst_n), .Q(x_z2[2])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[2]  ( .D(n1836), .CP(clk), .RN(rst_n), .Q(
        x_reg2[2]) );
  HS65_GS_DFPRQX4 \x_z2_reg[1]  ( .D(n1837), .CP(clk), .RN(rst_n), .Q(x_z2[1])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[1]  ( .D(n1838), .CP(clk), .RN(rst_n), .Q(
        x_reg2[1]) );
  HS65_GS_DFPRQX4 \x_z2_reg[0]  ( .D(n1839), .CP(clk), .RN(rst_n), .Q(x_z2[0])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[0]  ( .D(n1840), .CP(clk), .RN(rst_n), .Q(
        x_reg2[0]) );
  HS65_GS_DFPRQX4 \data_out_reg[15]  ( .D(n1841), .CP(clk), .RN(rst_n), .Q(
        data_out[15]) );
  HS65_GS_DFPRQX4 \y_z1_reg[15]  ( .D(n1842), .CP(clk), .RN(rst_n), .Q(
        y_z1[15]) );
  HS65_GS_DFPRQX4 \y_z2_reg[15]  ( .D(n1843), .CP(clk), .RN(rst_n), .Q(
        y_z2[15]) );
  HS65_GS_DFPRQX4 \data_out_reg[14]  ( .D(n1844), .CP(clk), .RN(rst_n), .Q(
        data_out[14]) );
  HS65_GS_DFPRQX4 \y_z1_reg[14]  ( .D(n1845), .CP(clk), .RN(rst_n), .Q(
        y_z1[14]) );
  HS65_GS_DFPRQX4 \y_z2_reg[14]  ( .D(n1846), .CP(clk), .RN(rst_n), .Q(
        y_z2[14]) );
  HS65_GS_DFPRQX4 \data_out_reg[13]  ( .D(n1847), .CP(clk), .RN(rst_n), .Q(
        data_out[13]) );
  HS65_GS_DFPRQX4 \y_z1_reg[13]  ( .D(n1848), .CP(clk), .RN(rst_n), .Q(
        y_z1[13]) );
  HS65_GS_DFPRQX4 \y_z2_reg[13]  ( .D(n1849), .CP(clk), .RN(rst_n), .Q(
        y_z2[13]) );
  HS65_GS_DFPRQX4 \data_out_reg[12]  ( .D(n1850), .CP(clk), .RN(rst_n), .Q(
        data_out[12]) );
  HS65_GS_DFPRQX4 \y_z1_reg[12]  ( .D(n1851), .CP(clk), .RN(rst_n), .Q(
        y_z1[12]) );
  HS65_GS_DFPRQX4 \y_z2_reg[12]  ( .D(n1852), .CP(clk), .RN(rst_n), .Q(
        y_z2[12]) );
  HS65_GS_DFPRQX4 \data_out_reg[11]  ( .D(n1853), .CP(clk), .RN(rst_n), .Q(
        data_out[11]) );
  HS65_GS_DFPRQX4 \y_z1_reg[11]  ( .D(n1854), .CP(clk), .RN(rst_n), .Q(
        y_z1[11]) );
  HS65_GS_DFPRQX4 \y_z2_reg[11]  ( .D(n1855), .CP(clk), .RN(rst_n), .Q(
        y_z2[11]) );
  HS65_GS_DFPRQX4 \data_out_reg[10]  ( .D(n1856), .CP(clk), .RN(rst_n), .Q(
        data_out[10]) );
  HS65_GS_DFPRQX4 \y_z1_reg[10]  ( .D(n1857), .CP(clk), .RN(rst_n), .Q(
        y_z1[10]) );
  HS65_GS_DFPRQX4 \y_z2_reg[10]  ( .D(n1858), .CP(clk), .RN(rst_n), .Q(
        y_z2[10]) );
  HS65_GS_DFPRQX4 \data_out_reg[9]  ( .D(n1859), .CP(clk), .RN(rst_n), .Q(
        data_out[9]) );
  HS65_GS_DFPRQX4 \y_z1_reg[9]  ( .D(n1860), .CP(clk), .RN(rst_n), .Q(y_z1[9])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[9]  ( .D(n1861), .CP(clk), .RN(rst_n), .Q(y_z2[9])
         );
  HS65_GS_DFPRQX4 \data_out_reg[8]  ( .D(n1862), .CP(clk), .RN(rst_n), .Q(
        data_out[8]) );
  HS65_GS_DFPRQX4 \y_z1_reg[8]  ( .D(n1863), .CP(clk), .RN(rst_n), .Q(y_z1[8])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[8]  ( .D(n1864), .CP(clk), .RN(rst_n), .Q(y_z2[8])
         );
  HS65_GS_DFPRQX4 \data_out_reg[7]  ( .D(n1865), .CP(clk), .RN(rst_n), .Q(
        data_out[7]) );
  HS65_GS_DFPRQX4 \y_z1_reg[7]  ( .D(n1866), .CP(clk), .RN(rst_n), .Q(y_z1[7])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[7]  ( .D(n1867), .CP(clk), .RN(rst_n), .Q(y_z2[7])
         );
  HS65_GS_DFPRQX4 \data_out_reg[6]  ( .D(n1868), .CP(clk), .RN(rst_n), .Q(
        data_out[6]) );
  HS65_GS_DFPRQX4 \y_z1_reg[6]  ( .D(n1869), .CP(clk), .RN(rst_n), .Q(y_z1[6])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[6]  ( .D(n1870), .CP(clk), .RN(rst_n), .Q(y_z2[6])
         );
  HS65_GS_DFPRQX4 \data_out_reg[5]  ( .D(n1871), .CP(clk), .RN(rst_n), .Q(
        data_out[5]) );
  HS65_GS_DFPRQX4 \y_z1_reg[5]  ( .D(n1872), .CP(clk), .RN(rst_n), .Q(y_z1[5])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[5]  ( .D(n1873), .CP(clk), .RN(rst_n), .Q(y_z2[5])
         );
  HS65_GS_DFPRQX4 \data_out_reg[4]  ( .D(n1874), .CP(clk), .RN(rst_n), .Q(
        data_out[4]) );
  HS65_GS_DFPRQX4 \y_z1_reg[4]  ( .D(n1875), .CP(clk), .RN(rst_n), .Q(y_z1[4])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[4]  ( .D(n1876), .CP(clk), .RN(rst_n), .Q(y_z2[4])
         );
  HS65_GS_DFPRQX4 \data_out_reg[3]  ( .D(n1877), .CP(clk), .RN(rst_n), .Q(
        data_out[3]) );
  HS65_GS_DFPRQX4 \y_z1_reg[3]  ( .D(n1878), .CP(clk), .RN(rst_n), .Q(y_z1[3])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[3]  ( .D(n1879), .CP(clk), .RN(rst_n), .Q(y_z2[3])
         );
  HS65_GS_DFPRQX4 \data_out_reg[2]  ( .D(n1880), .CP(clk), .RN(rst_n), .Q(
        data_out[2]) );
  HS65_GS_DFPRQX4 \y_z1_reg[2]  ( .D(n1881), .CP(clk), .RN(rst_n), .Q(y_z1[2])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[2]  ( .D(n1882), .CP(clk), .RN(rst_n), .Q(y_z2[2])
         );
  HS65_GS_DFPRQX4 \data_out_reg[1]  ( .D(n1883), .CP(clk), .RN(rst_n), .Q(
        data_out[1]) );
  HS65_GS_DFPRQX4 \y_z1_reg[1]  ( .D(n1884), .CP(clk), .RN(rst_n), .Q(y_z1[1])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[1]  ( .D(n1885), .CP(clk), .RN(rst_n), .Q(y_z2[1])
         );
  HS65_GS_DFPRQX4 \data_out_reg[0]  ( .D(n1886), .CP(clk), .RN(rst_n), .Q(
        data_out[0]) );
  HS65_GS_DFPRQX4 \y_z1_reg[0]  ( .D(n1887), .CP(clk), .RN(rst_n), .Q(y_z1[0])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[0]  ( .D(n1888), .CP(clk), .RN(rst_n), .Q(y_z2[0])
         );
  HS65_GS_IVX2 U3 ( .A(x_z2[15]), .Z(n1680) );
  HS65_GS_IVX2 U4 ( .A(x_z2[14]), .Z(n1682) );
  HS65_GS_IVX2 U5 ( .A(x_z2[13]), .Z(n1684) );
  HS65_GS_IVX2 U6 ( .A(x_z2[12]), .Z(n1686) );
  HS65_GS_IVX2 U7 ( .A(x_z2[11]), .Z(n1688) );
  HS65_GS_IVX2 U8 ( .A(x_z2[10]), .Z(n1690) );
  HS65_GS_IVX2 U9 ( .A(x_z2[9]), .Z(n1692) );
  HS65_GS_IVX2 U10 ( .A(x_z2[8]), .Z(n1694) );
  HS65_GS_IVX2 U11 ( .A(x_z2[7]), .Z(n1696) );
  HS65_GS_IVX2 U12 ( .A(x_z2[6]), .Z(n1698) );
  HS65_GS_IVX2 U13 ( .A(x_z2[5]), .Z(n1700) );
  HS65_GS_IVX2 U14 ( .A(x_z2[4]), .Z(n1702) );
  HS65_GS_IVX2 U15 ( .A(x_z2[3]), .Z(n1704) );
  HS65_GS_IVX2 U16 ( .A(x_z2[2]), .Z(n1706) );
  HS65_GS_HA1X4 U17 ( .A0(n1349), .B0(n1347), .CO(n1705) );
  HS65_GS_NOR2X3 U18 ( .A(x_z2[15]), .B(n1678), .Z(n1787) );
  HS65_GS_AND2X4 U19 ( .A(\mul_a2/fa1_c1_r[31] ), .B(\mul_a2/fa1_s2_r[32] ), 
        .Z(n139) );
  HS65_GS_AND2X4 U20 ( .A(\mul_a2/fa1_c1_r[30] ), .B(\mul_a2/fa1_s2_r[31] ), 
        .Z(n131) );
  HS65_GSS_XOR2X3 U21 ( .A(\mul_a2/fa1_s2_r[31] ), .B(\mul_a2/fa1_c1_r[30] ), 
        .Z(n128) );
  HS65_GS_AND2X4 U22 ( .A(n128), .B(\mul_a2/fa1_s0_r[31] ), .Z(n130) );
  HS65_GSS_XOR2X3 U23 ( .A(\mul_a2/fa1_s2_r[32] ), .B(\mul_a2/fa1_c1_r[31] ), 
        .Z(n1) );
  HS65_GSS_XOR2X3 U24 ( .A(n1), .B(\mul_a2/fa1_s0_r[32] ), .Z(n129) );
  HS65_GS_AND2X4 U25 ( .A(\mul_a2/fa1_s0_r[32] ), .B(n1), .Z(n2) );
  HS65_GSS_XOR2X3 U26 ( .A(n3), .B(n2), .Z(n136) );
  HS65_GS_FA1X4 U27 ( .A0(\mul_a2/fa1_c1_r[28] ), .B0(\mul_a2/fa1_c2_r[28] ), 
        .CI(\mul_a2/fa1_s2_r[29] ), .CO(n126), .S0(n4) );
  HS65_GS_AND2X4 U28 ( .A(\mul_a2/fa1_s0_r[29] ), .B(n4), .Z(n125) );
  HS65_GSS_XOR2X3 U29 ( .A(\mul_a2/fa1_s2_r[30] ), .B(\mul_a2/fa1_c1_r[29] ), 
        .Z(n127) );
  HS65_GSS_XOR2X3 U30 ( .A(\mul_a2/fa1_s0_r[30] ), .B(n127), .Z(n124) );
  HS65_GS_FA1X4 U31 ( .A0(\mul_a2/fa1_c1_r[27] ), .B0(\mul_a2/fa1_c2_r[27] ), 
        .CI(\mul_a2/fa1_s2_r[28] ), .CO(n123), .S0(n5) );
  HS65_GS_AND2X4 U32 ( .A(\mul_a2/fa1_s0_r[28] ), .B(n5), .Z(n122) );
  HS65_GSS_XOR2X3 U33 ( .A(n4), .B(\mul_a2/fa1_s0_r[29] ), .Z(n121) );
  HS65_GS_FA1X4 U34 ( .A0(\mul_a2/fa1_c1_r[26] ), .B0(\mul_a2/fa1_c2_r[26] ), 
        .CI(\mul_a2/fa1_s2_r[27] ), .CO(n120), .S0(n6) );
  HS65_GS_AND2X4 U35 ( .A(\mul_a2/fa1_s0_r[27] ), .B(n6), .Z(n119) );
  HS65_GSS_XOR2X3 U36 ( .A(n5), .B(\mul_a2/fa1_s0_r[28] ), .Z(n118) );
  HS65_GS_FA1X4 U37 ( .A0(\mul_a2/fa1_c1_r[25] ), .B0(\mul_a2/fa1_c2_r[25] ), 
        .CI(\mul_a2/fa1_s2_r[26] ), .CO(n117), .S0(n110) );
  HS65_GS_AND2X4 U38 ( .A(\mul_a2/fa1_s0_r[26] ), .B(n110), .Z(n116) );
  HS65_GSS_XOR2X3 U39 ( .A(n6), .B(\mul_a2/fa1_s0_r[27] ), .Z(n115) );
  HS65_GSS_XOR2X3 U40 ( .A(\mul_a2/fa1_s0_r[23] ), .B(\mul_a2/fa1_s1_r[23] ), 
        .Z(n98) );
  HS65_GS_FA1X4 U41 ( .A0(\mul_a2/fa1_c1_r[22] ), .B0(\mul_a2/fa1_c2_r[22] ), 
        .CI(\mul_a2/fa1_s2_r[23] ), .CO(n104), .S0(n97) );
  HS65_GS_AND2X4 U42 ( .A(\mul_a2/fa1_s0_r[22] ), .B(\mul_a2/fa1_s1_r[22] ), 
        .Z(n96) );
  HS65_GS_AND2X4 U43 ( .A(\mul_a2/fa1_s0_r[23] ), .B(\mul_a2/fa1_s1_r[23] ), 
        .Z(n105) );
  HS65_GS_FA1X4 U44 ( .A0(\mul_a2/fa1_c1_r[18] ), .B0(\mul_a2/fa1_c2_r[18] ), 
        .CI(\mul_a2/fa1_s2_r[19] ), .CO(n80), .S0(n9) );
  HS65_GSS_XOR2X3 U45 ( .A(\mul_a2/fa1_s0_r[19] ), .B(\mul_a2/fa1_s1_r[19] ), 
        .Z(n8) );
  HS65_GS_AND2X4 U46 ( .A(\mul_a2/fa1_s0_r[18] ), .B(\mul_a2/fa1_s1_r[18] ), 
        .Z(n7) );
  HS65_GS_AND2X4 U47 ( .A(\mul_a2/fa1_s0_r[19] ), .B(\mul_a2/fa1_s1_r[19] ), 
        .Z(n83) );
  HS65_GSS_XOR2X3 U48 ( .A(\mul_a2/fa1_s0_r[20] ), .B(\mul_a2/fa1_s1_r[20] ), 
        .Z(n81) );
  HS65_GS_FA1X4 U49 ( .A0(\mul_a2/fa1_c1_r[17] ), .B0(\mul_a2/fa1_c2_r[17] ), 
        .CI(\mul_a2/fa1_s2_r[18] ), .CO(n77), .S0(n12) );
  HS65_GSS_XOR2X3 U50 ( .A(\mul_a2/fa1_s0_r[18] ), .B(\mul_a2/fa1_s1_r[18] ), 
        .Z(n11) );
  HS65_GS_AND2X4 U51 ( .A(\mul_a2/fa1_s0_r[17] ), .B(\mul_a2/fa1_s1_r[17] ), 
        .Z(n10) );
  HS65_GS_FA1X4 U52 ( .A0(n9), .B0(n8), .CI(n7), .CO(n79), .S0(n75) );
  HS65_GS_FA1X4 U53 ( .A0(\mul_a2/fa1_c1_r[16] ), .B0(\mul_a2/fa1_c2_r[16] ), 
        .CI(\mul_a2/fa1_s2_r[17] ), .CO(n74), .S0(n15) );
  HS65_GSS_XOR2X3 U54 ( .A(\mul_a2/fa1_s0_r[17] ), .B(\mul_a2/fa1_s1_r[17] ), 
        .Z(n14) );
  HS65_GS_AND2X4 U55 ( .A(\mul_a2/fa1_s0_r[16] ), .B(\mul_a2/fa1_s1_r[16] ), 
        .Z(n13) );
  HS65_GS_FA1X4 U56 ( .A0(n12), .B0(n11), .CI(n10), .CO(n76), .S0(n72) );
  HS65_GSS_XOR2X3 U57 ( .A(\mul_a2/fa1_s0_r[16] ), .B(\mul_a2/fa1_s1_r[16] ), 
        .Z(n18) );
  HS65_GS_FA1X4 U58 ( .A0(\mul_a2/fa1_c1_r[15] ), .B0(\mul_a2/fa1_c2_r[15] ), 
        .CI(\mul_a2/fa1_s2_r[16] ), .CO(n71), .S0(n17) );
  HS65_GS_AND2X4 U59 ( .A(\mul_a2/fa1_s0_r[15] ), .B(\mul_a2/fa1_s1_r[15] ), 
        .Z(n16) );
  HS65_GS_FA1X4 U60 ( .A0(n15), .B0(n14), .CI(n13), .CO(n73), .S0(n69) );
  HS65_GS_FA1X4 U61 ( .A0(\mul_a2/fa1_c1_r[14] ), .B0(\mul_a2/fa1_c2_r[14] ), 
        .CI(\mul_a2/fa1_s2_r[15] ), .CO(n68), .S0(n21) );
  HS65_GSS_XOR2X3 U62 ( .A(\mul_a2/fa1_s0_r[15] ), .B(\mul_a2/fa1_s1_r[15] ), 
        .Z(n20) );
  HS65_GS_AND2X4 U63 ( .A(\mul_a2/fa1_s0_r[14] ), .B(\mul_a2/fa1_s1_r[14] ), 
        .Z(n19) );
  HS65_GS_FA1X4 U64 ( .A0(n18), .B0(n17), .CI(n16), .CO(n70), .S0(n66) );
  HS65_GS_AND2X4 U65 ( .A(\mul_a2/fa1_c1_r[13] ), .B(\mul_a2/fa1_s2_r[14] ), 
        .Z(n24) );
  HS65_GS_FA1X4 U66 ( .A0(n21), .B0(n20), .CI(n19), .CO(n67), .S0(n23) );
  HS65_GSS_XOR2X3 U67 ( .A(\mul_a2/fa1_c1_r[13] ), .B(\mul_a2/fa1_s2_r[14] ), 
        .Z(n62) );
  HS65_GSS_XOR2X3 U68 ( .A(\mul_a2/fa1_s0_r[14] ), .B(\mul_a2/fa1_s1_r[14] ), 
        .Z(n61) );
  HS65_GS_AND2X4 U69 ( .A(\mul_a2/fa1_s0_r[13] ), .B(\mul_a2/fa1_s1_r[13] ), 
        .Z(n60) );
  HS65_GS_FA1X4 U70 ( .A0(n24), .B0(n23), .CI(n22), .CO(n1607), .S0(n1611) );
  HS65_GSS_XOR2X3 U71 ( .A(\mul_a2/fa1_s0_r[11] ), .B(\mul_a2/fa1_s1_r[11] ), 
        .Z(n31) );
  HS65_GS_AND2X4 U72 ( .A(\mul_a2/fa1_s0_r[10] ), .B(\mul_a2/fa1_s1_r[10] ), 
        .Z(n30) );
  HS65_GSS_XOR2X3 U73 ( .A(\mul_a2/fa1_s2_r[12] ), .B(\mul_a2/fa1_c1_r[11] ), 
        .Z(n27) );
  HS65_GSS_XOR2X3 U74 ( .A(\mul_a2/fa1_s0_r[12] ), .B(\mul_a2/fa1_s1_r[12] ), 
        .Z(n26) );
  HS65_GS_AND2X4 U75 ( .A(\mul_a2/fa1_s0_r[11] ), .B(\mul_a2/fa1_s1_r[11] ), 
        .Z(n25) );
  HS65_GS_AND2X4 U76 ( .A(n28), .B(n29), .Z(n53) );
  HS65_GS_AND2X4 U77 ( .A(\mul_a2/fa1_s2_r[12] ), .B(\mul_a2/fa1_c1_r[11] ), 
        .Z(n56) );
  HS65_GS_FA1X4 U78 ( .A0(n27), .B0(n26), .CI(n25), .CO(n55), .S0(n29) );
  HS65_GS_AND2X4 U79 ( .A(\mul_a2/fa1_s0_r[12] ), .B(\mul_a2/fa1_s1_r[12] ), 
        .Z(n59) );
  HS65_GSS_XOR2X3 U80 ( .A(\mul_a2/fa1_s2_r[13] ), .B(\mul_a2/fa1_c1_r[12] ), 
        .Z(n58) );
  HS65_GSS_XOR2X3 U81 ( .A(\mul_a2/fa1_s0_r[13] ), .B(\mul_a2/fa1_s1_r[13] ), 
        .Z(n57) );
  HS65_GSS_XOR2X3 U82 ( .A(n29), .B(n28), .Z(n50) );
  HS65_GS_AND2X4 U83 ( .A(\mul_a2/fa1_s0_r[9] ), .B(\mul_a2/fa1_s1_r[9] ), .Z(
        n37) );
  HS65_GSS_XOR2X3 U84 ( .A(\mul_a2/fa1_s0_r[10] ), .B(\mul_a2/fa1_s1_r[10] ), 
        .Z(n36) );
  HS65_GS_FA1X4 U85 ( .A0(\mul_a2/fa1_c1_r[10] ), .B0(n31), .CI(n30), .CO(n28), 
        .S0(n44) );
  HS65_GS_AND2X4 U86 ( .A(n43), .B(n44), .Z(n49) );
  HS65_GSS_XOR2X3 U87 ( .A(\mul_a2/fa1_s0_r[9] ), .B(\mul_a2/fa1_s1_r[9] ), 
        .Z(n40) );
  HS65_GS_AND2X4 U88 ( .A(\mul_a2/fa1_s0_r[8] ), .B(\mul_a2/fa1_s1_r[8] ), .Z(
        n39) );
  HS65_GS_AND2X4 U89 ( .A(\mul_a2/fa1_s0_r[7] ), .B(\mul_a2/fa1_s1_r[7] ), .Z(
        n33) );
  HS65_GSS_XOR2X3 U90 ( .A(\mul_a2/fa1_s0_r[8] ), .B(\mul_a2/fa1_s1_r[8] ), 
        .Z(n32) );
  HS65_GS_AND2X4 U91 ( .A(n33), .B(n32), .Z(n34) );
  HS65_GS_AND2X4 U92 ( .A(n35), .B(n34), .Z(n38) );
  HS65_GS_FA1X4 U93 ( .A0(n37), .B0(\mul_a2/fa1_c1_r[9] ), .CI(n36), .CO(n43), 
        .S0(n41) );
  HS65_GS_AND2X4 U94 ( .A(n38), .B(n41), .Z(n47) );
  HS65_GS_FA1X4 U95 ( .A0(\mul_a2/fa1_c1_r[8] ), .B0(n40), .CI(n39), .CO(n42), 
        .S0(n35) );
  HS65_GS_AND2X4 U96 ( .A(n42), .B(n41), .Z(n46) );
  HS65_GSS_XOR2X3 U97 ( .A(n44), .B(n43), .Z(n45) );
  HS65_GS_PAO2X4 U98 ( .A(n47), .B(n46), .P(n45), .Z(n48) );
  HS65_GS_PAO2X4 U99 ( .A(n50), .B(n49), .P(n48), .Z(n51) );
  HS65_GS_PAO2X4 U100 ( .A(n53), .B(n52), .P(n51), .Z(n1615) );
  HS65_GS_FA1X4 U101 ( .A0(n56), .B0(n55), .CI(n54), .CO(n1614), .S0(n52) );
  HS65_GS_FA1X4 U102 ( .A0(n59), .B0(n58), .CI(n57), .CO(n65), .S0(n54) );
  HS65_GS_AND2X4 U103 ( .A(\mul_a2/fa1_s2_r[13] ), .B(\mul_a2/fa1_c1_r[12] ), 
        .Z(n64) );
  HS65_GS_FA1X4 U104 ( .A0(n62), .B0(n61), .CI(n60), .CO(n22), .S0(n63) );
  HS65_GS_FA1X4 U105 ( .A0(n65), .B0(n64), .CI(n63), .CO(n1609), .S0(n1613) );
  HS65_GS_FA1X4 U106 ( .A0(n68), .B0(n67), .CI(n66), .CO(n1603), .S0(n1605) );
  HS65_GS_FA1X4 U107 ( .A0(n71), .B0(n70), .CI(n69), .CO(n1599), .S0(n1601) );
  HS65_GS_FA1X4 U108 ( .A0(n74), .B0(n73), .CI(n72), .CO(n1595), .S0(n1597) );
  HS65_GS_FA1X4 U109 ( .A0(n77), .B0(n76), .CI(n75), .CO(n1591), .S0(n1593) );
  HS65_GS_FA1X4 U110 ( .A0(n80), .B0(n79), .CI(n78), .CO(n1587), .S0(n1589) );
  HS65_GS_FA1X4 U111 ( .A0(\mul_a2/fa1_c1_r[19] ), .B0(\mul_a2/fa1_c2_r[19] ), 
        .CI(\mul_a2/fa1_s2_r[20] ), .CO(n86), .S0(n82) );
  HS65_GS_FA1X4 U112 ( .A0(n83), .B0(n82), .CI(n81), .CO(n85), .S0(n78) );
  HS65_GSS_XOR2X3 U113 ( .A(\mul_a2/fa1_s0_r[21] ), .B(\mul_a2/fa1_s1_r[21] ), 
        .Z(n88) );
  HS65_GS_AND2X4 U114 ( .A(\mul_a2/fa1_s0_r[20] ), .B(\mul_a2/fa1_s1_r[20] ), 
        .Z(n87) );
  HS65_GS_FA1X4 U115 ( .A0(n86), .B0(n85), .CI(n84), .CO(n1582), .S0(n1585) );
  HS65_GS_FA1X4 U116 ( .A0(\mul_a2/fa1_c1_r[20] ), .B0(\mul_a2/fa1_c2_r[20] ), 
        .CI(\mul_a2/fa1_s2_r[21] ), .CO(n92), .S0(n89) );
  HS65_GS_FA1X4 U117 ( .A0(n89), .B0(n88), .CI(n87), .CO(n91), .S0(n84) );
  HS65_GS_AND2X4 U118 ( .A(\mul_a2/fa1_s0_r[21] ), .B(\mul_a2/fa1_s1_r[21] ), 
        .Z(n95) );
  HS65_GSS_XOR2X3 U119 ( .A(\mul_a2/fa1_s0_r[22] ), .B(\mul_a2/fa1_s1_r[22] ), 
        .Z(n93) );
  HS65_GS_FA1X4 U120 ( .A0(n92), .B0(n91), .CI(n90), .CO(n1578), .S0(n1581) );
  HS65_GS_FA1X4 U121 ( .A0(\mul_a2/fa1_c1_r[21] ), .B0(\mul_a2/fa1_c2_r[21] ), 
        .CI(\mul_a2/fa1_s2_r[22] ), .CO(n101), .S0(n94) );
  HS65_GS_FA1X4 U122 ( .A0(n95), .B0(n94), .CI(n93), .CO(n100), .S0(n90) );
  HS65_GS_FA1X4 U123 ( .A0(n98), .B0(n97), .CI(n96), .CO(n103), .S0(n99) );
  HS65_GS_FA1X4 U124 ( .A0(n101), .B0(n100), .CI(n99), .CO(n1574), .S0(n1577)
         );
  HS65_GS_FA1X4 U125 ( .A0(n104), .B0(n103), .CI(n102), .CO(n1571), .S0(n1573)
         );
  HS65_GS_FA1X4 U126 ( .A0(\mul_a2/fa1_c1_r[23] ), .B0(\mul_a2/fa1_c2_r[23] ), 
        .CI(\mul_a2/fa1_s2_r[24] ), .CO(n109), .S0(n106) );
  HS65_GS_FA1X4 U127 ( .A0(n106), .B0(\mul_a2/fa1_s0_r[24] ), .CI(n105), .CO(
        n108), .S0(n102) );
  HS65_GSS_XOR2X3 U128 ( .A(\mul_a2/fa1_s0_r[25] ), .B(n111), .Z(n107) );
  HS65_GS_FA1X4 U129 ( .A0(n109), .B0(n108), .CI(n107), .CO(n1566), .S0(n1569)
         );
  HS65_GSS_XOR2X3 U130 ( .A(n110), .B(\mul_a2/fa1_s0_r[26] ), .Z(n114) );
  HS65_GS_FA1X4 U131 ( .A0(\mul_a2/fa1_c1_r[24] ), .B0(\mul_a2/fa1_c2_r[24] ), 
        .CI(\mul_a2/fa1_s2_r[25] ), .CO(n113), .S0(n111) );
  HS65_GS_AND2X4 U132 ( .A(n111), .B(\mul_a2/fa1_s0_r[25] ), .Z(n112) );
  HS65_GS_FA1X4 U133 ( .A0(n114), .B0(n113), .CI(n112), .CO(n1562), .S0(n1565)
         );
  HS65_GS_FA1X4 U134 ( .A0(n117), .B0(n116), .CI(n115), .CO(n1540), .S0(n1561)
         );
  HS65_GS_FA1X4 U135 ( .A0(n120), .B0(n119), .CI(n118), .CO(n1550), .S0(n1538)
         );
  HS65_GS_FA1X4 U136 ( .A0(n123), .B0(n122), .CI(n121), .CO(n1547), .S0(n1548)
         );
  HS65_GS_FA1X4 U137 ( .A0(n126), .B0(n125), .CI(n124), .CO(n1543), .S0(n1545)
         );
  HS65_GS_AND2X4 U138 ( .A(\mul_a2/fa1_c1_r[29] ), .B(\mul_a2/fa1_s2_r[30] ), 
        .Z(n134) );
  HS65_GS_AND2X4 U139 ( .A(n127), .B(\mul_a2/fa1_s0_r[30] ), .Z(n133) );
  HS65_GSS_XOR2X3 U140 ( .A(\mul_a2/fa1_s0_r[31] ), .B(n128), .Z(n132) );
  HS65_GS_FA1X4 U141 ( .A0(n131), .B0(n130), .CI(n129), .CO(n3), .S0(n1552) );
  HS65_GS_FA1X4 U142 ( .A0(n134), .B0(n133), .CI(n132), .CO(n1551), .S0(n1541)
         );
  HS65_GSS_XOR2X3 U143 ( .A(n136), .B(n135), .Z(n137) );
  HS65_GSS_XOR3X2 U144 ( .A(\mul_a2/fa1_s0_r[33] ), .B(\mul_a2/fa1_c1_r[32] ), 
        .C(n137), .Z(n138) );
  HS65_GSS_XOR3X2 U145 ( .A(n139), .B(\mul_a2/fa1_s2_r[33] ), .C(n138), .Z(
        \mul_a2/result_sat[15] ) );
  HS65_GS_AND2X4 U146 ( .A(\mul_b2/fa1_s1_r[31] ), .B(\mul_b2/fa1_c0_r[30] ), 
        .Z(n233) );
  HS65_GSS_XOR2X3 U147 ( .A(\mul_b2/fa1_s1_r[32] ), .B(\mul_b2/fa1_c0_r[31] ), 
        .Z(n232) );
  HS65_GS_AND2X4 U148 ( .A(\mul_b2/fa1_s1_r[30] ), .B(\mul_b2/fa1_c0_r[29] ), 
        .Z(n141) );
  HS65_GSS_XOR2X3 U149 ( .A(\mul_b2/fa1_s1_r[31] ), .B(\mul_b2/fa1_c0_r[30] ), 
        .Z(n140) );
  HS65_GS_FA1X4 U150 ( .A0(\mul_b2/fa1_s2_r[31] ), .B0(n141), .CI(n140), .CO(
        n823), .S0(n815) );
  HS65_GS_AND2X4 U151 ( .A(\mul_b2/fa1_c0_r[28] ), .B(\mul_b2/fa1_s1_r[29] ), 
        .Z(n143) );
  HS65_GSS_XOR2X3 U152 ( .A(\mul_b2/fa1_s1_r[30] ), .B(\mul_b2/fa1_c0_r[29] ), 
        .Z(n142) );
  HS65_GS_FA1X4 U153 ( .A0(\mul_b2/fa1_s2_r[30] ), .B0(n143), .CI(n142), .CO(
        n814), .S0(n818) );
  HS65_GS_AND2X4 U154 ( .A(\mul_b2/fa1_c0_r[27] ), .B(\mul_b2/fa1_s1_r[28] ), 
        .Z(n145) );
  HS65_GSS_XOR2X3 U155 ( .A(\mul_b2/fa1_c0_r[28] ), .B(\mul_b2/fa1_s1_r[29] ), 
        .Z(n144) );
  HS65_GS_FA1X4 U156 ( .A0(\mul_b2/fa1_s2_r[29] ), .B0(n145), .CI(n144), .CO(
        n817), .S0(n821) );
  HS65_GS_AND2X4 U157 ( .A(\mul_b2/fa1_c0_r[26] ), .B(\mul_b2/fa1_s1_r[27] ), 
        .Z(n147) );
  HS65_GSS_XOR2X3 U158 ( .A(\mul_b2/fa1_c0_r[27] ), .B(\mul_b2/fa1_s1_r[28] ), 
        .Z(n146) );
  HS65_GS_FA1X4 U159 ( .A0(\mul_b2/fa1_s2_r[28] ), .B0(n147), .CI(n146), .CO(
        n820), .S0(n1012) );
  HS65_GS_AND2X4 U160 ( .A(\mul_b2/fa1_c0_r[25] ), .B(\mul_b2/fa1_s1_r[26] ), 
        .Z(n149) );
  HS65_GSS_XOR2X3 U161 ( .A(\mul_b2/fa1_c0_r[26] ), .B(\mul_b2/fa1_s1_r[27] ), 
        .Z(n148) );
  HS65_GS_FA1X4 U162 ( .A0(\mul_b2/fa1_s2_r[27] ), .B0(n149), .CI(n148), .CO(
        n1011), .S0(n1016) );
  HS65_GS_AND2X4 U163 ( .A(\mul_b2/fa1_c0_r[24] ), .B(\mul_b2/fa1_s1_r[25] ), 
        .Z(n226) );
  HS65_GSS_XOR2X3 U164 ( .A(\mul_b2/fa1_c0_r[25] ), .B(\mul_b2/fa1_s1_r[26] ), 
        .Z(n225) );
  HS65_GS_AND2X4 U165 ( .A(\mul_b2/fa1_c0_r[22] ), .B(\mul_b2/fa1_s1_r[23] ), 
        .Z(n151) );
  HS65_GSS_XOR2X3 U166 ( .A(\mul_b2/fa1_s1_r[24] ), .B(\mul_b2/fa1_c0_r[23] ), 
        .Z(n150) );
  HS65_GS_AND2X4 U167 ( .A(\mul_b2/fa1_s1_r[24] ), .B(\mul_b2/fa1_c0_r[23] ), 
        .Z(n228) );
  HS65_GSS_XOR2X3 U168 ( .A(\mul_b2/fa1_c0_r[24] ), .B(\mul_b2/fa1_s1_r[25] ), 
        .Z(n227) );
  HS65_GS_AND2X4 U169 ( .A(\mul_b2/fa1_c0_r[21] ), .B(\mul_b2/fa1_s1_r[22] ), 
        .Z(n153) );
  HS65_GSS_XOR2X3 U170 ( .A(\mul_b2/fa1_c0_r[22] ), .B(\mul_b2/fa1_s1_r[23] ), 
        .Z(n152) );
  HS65_GS_FA1X4 U171 ( .A0(\mul_b2/fa1_s2_r[24] ), .B0(n151), .CI(n150), .CO(
        n224), .S0(n220) );
  HS65_GS_AND2X4 U172 ( .A(\mul_b2/fa1_c0_r[20] ), .B(\mul_b2/fa1_s1_r[21] ), 
        .Z(n155) );
  HS65_GSS_XOR2X3 U173 ( .A(\mul_b2/fa1_c0_r[21] ), .B(\mul_b2/fa1_s1_r[22] ), 
        .Z(n154) );
  HS65_GS_FA1X4 U174 ( .A0(\mul_b2/fa1_s2_r[23] ), .B0(n153), .CI(n152), .CO(
        n221), .S0(n217) );
  HS65_GS_AND2X4 U175 ( .A(\mul_b2/fa1_c0_r[19] ), .B(\mul_b2/fa1_s1_r[20] ), 
        .Z(n157) );
  HS65_GSS_XOR2X3 U176 ( .A(\mul_b2/fa1_c0_r[20] ), .B(\mul_b2/fa1_s1_r[21] ), 
        .Z(n156) );
  HS65_GS_FA1X4 U177 ( .A0(\mul_b2/fa1_s2_r[22] ), .B0(n155), .CI(n154), .CO(
        n218), .S0(n214) );
  HS65_GS_AND2X4 U178 ( .A(\mul_b2/fa1_c0_r[18] ), .B(\mul_b2/fa1_s1_r[19] ), 
        .Z(n159) );
  HS65_GSS_XOR2X3 U179 ( .A(\mul_b2/fa1_c0_r[19] ), .B(\mul_b2/fa1_s1_r[20] ), 
        .Z(n158) );
  HS65_GS_FA1X4 U180 ( .A0(\mul_b2/fa1_s2_r[21] ), .B0(n157), .CI(n156), .CO(
        n215), .S0(n211) );
  HS65_GS_PAO2X4 U181 ( .A(\mul_b2/fa1_s1_r[18] ), .B(\mul_b2/fa1_s0_r[18] ), 
        .P(\mul_b2/fa1_c0_r[17] ), .Z(n161) );
  HS65_GSS_XOR2X3 U182 ( .A(\mul_b2/fa1_c0_r[18] ), .B(\mul_b2/fa1_s1_r[19] ), 
        .Z(n160) );
  HS65_GS_FA1X4 U183 ( .A0(\mul_b2/fa1_s2_r[20] ), .B0(n159), .CI(n158), .CO(
        n212), .S0(n208) );
  HS65_GS_FA1X4 U184 ( .A0(\mul_b2/fa1_s2_r[19] ), .B0(n161), .CI(n160), .CO(
        n209), .S0(n857) );
  HS65_GSS_XOR3X2 U185 ( .A(\mul_b2/fa1_s1_r[18] ), .B(\mul_b2/fa1_s0_r[18] ), 
        .C(\mul_b2/fa1_c0_r[17] ), .Z(n206) );
  HS65_GS_PAO2X4 U186 ( .A(\mul_b2/fa1_c0_r[16] ), .B(\mul_b2/fa1_s1_r[17] ), 
        .P(\mul_b2/fa1_s0_r[17] ), .Z(n205) );
  HS65_GS_PAO2X4 U187 ( .A(\mul_b2/fa1_s1_r[15] ), .B(\mul_b2/fa1_s0_r[15] ), 
        .P(\mul_b2/fa1_c0_r[14] ), .Z(n163) );
  HS65_GSS_XOR3X2 U188 ( .A(\mul_b2/fa1_c0_r[15] ), .B(\mul_b2/fa1_s1_r[16] ), 
        .C(\mul_b2/fa1_s0_r[16] ), .Z(n162) );
  HS65_GS_PAO2X4 U189 ( .A(\mul_b2/fa1_c0_r[15] ), .B(\mul_b2/fa1_s1_r[16] ), 
        .P(\mul_b2/fa1_s0_r[16] ), .Z(n204) );
  HS65_GSS_XOR3X2 U190 ( .A(\mul_b2/fa1_c0_r[16] ), .B(\mul_b2/fa1_s1_r[17] ), 
        .C(\mul_b2/fa1_s0_r[17] ), .Z(n203) );
  HS65_GSS_XOR3X2 U191 ( .A(\mul_b2/fa1_s1_r[15] ), .B(\mul_b2/fa1_s0_r[15] ), 
        .C(\mul_b2/fa1_c0_r[14] ), .Z(n165) );
  HS65_GS_PAO2X4 U192 ( .A(\mul_b2/fa1_s1_r[14] ), .B(\mul_b2/fa1_s0_r[14] ), 
        .P(\mul_b2/fa1_c0_r[13] ), .Z(n164) );
  HS65_GS_FA1X4 U193 ( .A0(\mul_b2/fa1_s2_r[16] ), .B0(n163), .CI(n162), .CO(
        n1028), .S0(n1031) );
  HS65_GS_FA1X4 U194 ( .A0(\mul_b2/fa1_s2_r[15] ), .B0(n165), .CI(n164), .CO(
        n1032), .S0(n167) );
  HS65_GSS_XOR3X2 U195 ( .A(\mul_b2/fa1_s1_r[14] ), .B(\mul_b2/fa1_s0_r[14] ), 
        .C(\mul_b2/fa1_c0_r[13] ), .Z(n169) );
  HS65_GS_PAO2X4 U196 ( .A(\mul_b2/fa1_s1_r[13] ), .B(\mul_b2/fa1_s0_r[13] ), 
        .P(\mul_b2/fa1_c0_r[12] ), .Z(n168) );
  HS65_GS_NOR2X2 U197 ( .A(n166), .B(n167), .Z(n202) );
  HS65_GS_AOI12X2 U198 ( .A(n167), .B(n166), .C(n202), .Z(n863) );
  HS65_GS_PAO2X4 U199 ( .A(\mul_b2/fa1_s1_r[12] ), .B(\mul_b2/fa1_s0_r[12] ), 
        .P(\mul_b2/fa1_c0_r[11] ), .Z(n171) );
  HS65_GSS_XOR3X2 U200 ( .A(\mul_b2/fa1_s1_r[13] ), .B(\mul_b2/fa1_s0_r[13] ), 
        .C(\mul_b2/fa1_c0_r[12] ), .Z(n170) );
  HS65_GS_FA1X4 U201 ( .A0(\mul_b2/fa1_s2_r[14] ), .B0(n169), .CI(n168), .CO(
        n166), .S0(n200) );
  HS65_GS_FA1X4 U202 ( .A0(\mul_b2/fa1_s2_r[13] ), .B0(n171), .CI(n170), .CO(
        n201), .S0(n198) );
  HS65_GSS_XOR3X2 U203 ( .A(\mul_b2/fa1_s1_r[12] ), .B(\mul_b2/fa1_s0_r[12] ), 
        .C(\mul_b2/fa1_c0_r[11] ), .Z(n191) );
  HS65_GS_PAO2X4 U204 ( .A(\mul_b2/fa1_c0_r[10] ), .B(\mul_b2/fa1_s1_r[11] ), 
        .P(\mul_b2/fa1_s0_r[11] ), .Z(n190) );
  HS65_GSS_XOR3X2 U205 ( .A(\mul_b2/fa1_c0_r[10] ), .B(\mul_b2/fa1_s1_r[11] ), 
        .C(\mul_b2/fa1_s0_r[11] ), .Z(n195) );
  HS65_GS_PAO2X4 U206 ( .A(\mul_b2/fa1_c0_r[9] ), .B(\mul_b2/fa1_s1_r[10] ), 
        .P(\mul_b2/fa1_s0_r[10] ), .Z(n194) );
  HS65_GS_PAO2X4 U207 ( .A(\mul_b2/fa1_s1_r[9] ), .B(\mul_b2/fa1_s0_r[9] ), 
        .P(\mul_b2/fa1_c0_r[8] ), .Z(n185) );
  HS65_GSS_XOR3X2 U208 ( .A(\mul_b2/fa1_c0_r[9] ), .B(\mul_b2/fa1_s1_r[10] ), 
        .C(\mul_b2/fa1_s0_r[10] ), .Z(n184) );
  HS65_GS_NOR2X2 U209 ( .A(n185), .B(n184), .Z(n189) );
  HS65_GS_PAO2X4 U210 ( .A(\mul_b2/fa1_c0_r[7] ), .B(\mul_b2/fa1_s1_r[8] ), 
        .P(\mul_b2/fa1_s0_r[8] ), .Z(n182) );
  HS65_GSS_XOR3X2 U211 ( .A(\mul_b2/fa1_s1_r[9] ), .B(\mul_b2/fa1_s0_r[9] ), 
        .C(\mul_b2/fa1_c0_r[8] ), .Z(n181) );
  HS65_GS_PAO2X4 U212 ( .A(\mul_b2/fa1_c0_r[5] ), .B(\mul_b2/fa1_s1_r[6] ), 
        .P(\mul_b2/fa1_s0_r[6] ), .Z(n176) );
  HS65_GSS_XOR3X2 U213 ( .A(\mul_b2/fa1_c0_r[6] ), .B(\mul_b2/fa1_s1_r[7] ), 
        .C(\mul_b2/fa1_s0_r[7] ), .Z(n175) );
  HS65_GS_NAND2X2 U214 ( .A(\mul_b2/fa1_s0_r[5] ), .B(\mul_b2/fa1_c0_r[4] ), 
        .Z(n173) );
  HS65_GSS_XNOR3X2 U215 ( .A(\mul_b2/fa1_c0_r[5] ), .B(\mul_b2/fa1_s1_r[6] ), 
        .C(\mul_b2/fa1_s0_r[6] ), .Z(n172) );
  HS65_GS_NOR2X2 U216 ( .A(n173), .B(n172), .Z(n174) );
  HS65_GS_PAO2X4 U217 ( .A(n176), .B(n175), .P(n174), .Z(n179) );
  HS65_GS_PAO2X4 U218 ( .A(\mul_b2/fa1_c0_r[6] ), .B(\mul_b2/fa1_s1_r[7] ), 
        .P(\mul_b2/fa1_s0_r[7] ), .Z(n178) );
  HS65_GSS_XOR3X2 U219 ( .A(\mul_b2/fa1_c0_r[7] ), .B(\mul_b2/fa1_s1_r[8] ), 
        .C(\mul_b2/fa1_s0_r[8] ), .Z(n177) );
  HS65_GS_PAO2X4 U220 ( .A(n179), .B(n178), .P(n177), .Z(n180) );
  HS65_GS_OAI21X2 U221 ( .A(n182), .B(n181), .C(n180), .Z(n188) );
  HS65_GS_AND2X4 U222 ( .A(n182), .B(n181), .Z(n183) );
  HS65_GS_PAOI2X1 U223 ( .A(n185), .B(n184), .P(n183), .Z(n187) );
  HS65_GS_NOR2X2 U224 ( .A(n194), .B(n195), .Z(n186) );
  HS65_GS_CBI4I6X2 U225 ( .A(n189), .B(n188), .C(n187), .D(n186), .Z(n193) );
  HS65_GS_FA1X4 U226 ( .A0(\mul_b2/fa1_s2_r[12] ), .B0(n191), .CI(n190), .CO(
        n197), .S0(n192) );
  HS65_GS_CB4I1X4 U227 ( .A(n195), .B(n194), .C(n193), .D(n192), .Z(n196) );
  HS65_GS_PAOI2X1 U228 ( .A(n198), .B(n197), .P(n196), .Z(n866) );
  HS65_GS_NAND2X2 U229 ( .A(n200), .B(n201), .Z(n199) );
  HS65_GS_OAI21X2 U230 ( .A(n200), .B(n201), .C(n199), .Z(n865) );
  HS65_GS_NOR2X2 U231 ( .A(n866), .B(n865), .Z(n864) );
  HS65_GS_AOI12X2 U232 ( .A(n201), .B(n200), .C(n864), .Z(n862) );
  HS65_GS_AOI12X2 U233 ( .A(n863), .B(n862), .C(n202), .Z(n1030) );
  HS65_GS_FA1X4 U234 ( .A0(\mul_b2/fa1_s2_r[17] ), .B0(n204), .CI(n203), .CO(
        n1023), .S0(n1027) );
  HS65_GS_FA1X4 U235 ( .A0(\mul_b2/fa1_s2_r[18] ), .B0(n206), .CI(n205), .CO(
        n856), .S0(n1022) );
  HS65_GS_PAOI2X1 U236 ( .A(n857), .B(n856), .P(n859), .Z(n854) );
  HS65_GS_NAND2X2 U237 ( .A(n208), .B(n209), .Z(n207) );
  HS65_GS_OAI21X2 U238 ( .A(n208), .B(n209), .C(n207), .Z(n853) );
  HS65_GS_NOR2X2 U239 ( .A(n854), .B(n853), .Z(n852) );
  HS65_GS_AOI12X2 U240 ( .A(n209), .B(n208), .C(n852), .Z(n850) );
  HS65_GS_NAND2X2 U241 ( .A(n211), .B(n212), .Z(n210) );
  HS65_GS_OAI21X2 U242 ( .A(n211), .B(n212), .C(n210), .Z(n849) );
  HS65_GS_NOR2X2 U243 ( .A(n850), .B(n849), .Z(n848) );
  HS65_GS_AOI12X2 U244 ( .A(n212), .B(n211), .C(n848), .Z(n846) );
  HS65_GS_NAND2X2 U245 ( .A(n214), .B(n215), .Z(n213) );
  HS65_GS_OAI21X2 U246 ( .A(n214), .B(n215), .C(n213), .Z(n845) );
  HS65_GS_NOR2X2 U247 ( .A(n846), .B(n845), .Z(n844) );
  HS65_GS_AOI12X2 U248 ( .A(n215), .B(n214), .C(n844), .Z(n842) );
  HS65_GS_NAND2X2 U249 ( .A(n217), .B(n218), .Z(n216) );
  HS65_GS_OAI21X2 U250 ( .A(n217), .B(n218), .C(n216), .Z(n841) );
  HS65_GS_NOR2X2 U251 ( .A(n842), .B(n841), .Z(n840) );
  HS65_GS_AOI12X2 U252 ( .A(n218), .B(n217), .C(n840), .Z(n838) );
  HS65_GS_NAND2X2 U253 ( .A(n220), .B(n221), .Z(n219) );
  HS65_GS_OAI21X2 U254 ( .A(n220), .B(n221), .C(n219), .Z(n837) );
  HS65_GS_NOR2X2 U255 ( .A(n838), .B(n837), .Z(n836) );
  HS65_GS_AOI12X2 U256 ( .A(n221), .B(n220), .C(n836), .Z(n834) );
  HS65_GS_NAND2X2 U257 ( .A(n223), .B(n224), .Z(n222) );
  HS65_GS_OAI21X2 U258 ( .A(n223), .B(n224), .C(n222), .Z(n833) );
  HS65_GS_NOR2X2 U259 ( .A(n834), .B(n833), .Z(n832) );
  HS65_GS_AOI12X2 U260 ( .A(n224), .B(n223), .C(n832), .Z(n1020) );
  HS65_GS_FA1X4 U261 ( .A0(\mul_b2/fa1_s2_r[26] ), .B0(n226), .CI(n225), .CO(
        n1015), .S0(n230) );
  HS65_GS_FA1X4 U262 ( .A0(\mul_b2/fa1_s2_r[25] ), .B0(n228), .CI(n227), .CO(
        n229), .S0(n223) );
  HS65_GS_NAND2X2 U263 ( .A(n230), .B(n229), .Z(n231) );
  HS65_GS_OAI21X2 U264 ( .A(n230), .B(n229), .C(n231), .Z(n1021) );
  HS65_GS_OAI21X2 U265 ( .A(n1020), .B(n1021), .C(n231), .Z(n1014) );
  HS65_GS_NAND2X2 U266 ( .A(\mul_b2/fa1_s1_r[32] ), .B(\mul_b2/fa1_c0_r[31] ), 
        .Z(n235) );
  HS65_GS_FA1X4 U267 ( .A0(\mul_b2/fa1_s2_r[32] ), .B0(n233), .CI(n232), .CO(
        n234), .S0(n824) );
  HS65_GSS_XNOR2X3 U268 ( .A(n235), .B(n234), .Z(n236) );
  HS65_GSS_XOR3X2 U269 ( .A(\mul_b2/fa1_c0_r[32] ), .B(n237), .C(n236), .Z(
        n238) );
  HS65_GSS_XOR3X2 U270 ( .A(n238), .B(\mul_b2/fa1_s1_r[33] ), .C(
        \mul_b2/fa1_s2_r[33] ), .Z(\mul_b2/result_sat[15] ) );
  HS65_GSS_XOR2X3 U271 ( .A(\mul_b0/fa1_s0_r[32] ), .B(\mul_b0/fa1_s1_r[32] ), 
        .Z(n240) );
  HS65_GS_AND2X4 U272 ( .A(\mul_b0/fa1_s0_r[31] ), .B(\mul_b0/fa1_s1_r[31] ), 
        .Z(n239) );
  HS65_GS_AND2X4 U273 ( .A(\mul_b0/fa1_s1_r[32] ), .B(\mul_b0/fa1_s0_r[32] ), 
        .Z(n352) );
  HS65_GSS_XOR2X3 U274 ( .A(\mul_b0/fa1_s0_r[30] ), .B(\mul_b0/fa1_s1_r[30] ), 
        .Z(n244) );
  HS65_GS_AND2X4 U275 ( .A(\mul_b0/fa1_s0_r[29] ), .B(\mul_b0/fa1_s1_r[29] ), 
        .Z(n243) );
  HS65_GSS_XOR2X3 U276 ( .A(\mul_b0/fa1_s0_r[31] ), .B(\mul_b0/fa1_s1_r[31] ), 
        .Z(n242) );
  HS65_GS_AND2X4 U277 ( .A(\mul_b0/fa1_s0_r[30] ), .B(\mul_b0/fa1_s1_r[30] ), 
        .Z(n241) );
  HS65_GS_FA1X4 U278 ( .A0(\mul_b0/fa1_s2_r[32] ), .B0(n240), .CI(n239), .CO(
        n353), .S0(n349) );
  HS65_GS_FA1X4 U279 ( .A0(\mul_b0/fa1_s2_r[31] ), .B0(n242), .CI(n241), .CO(
        n348), .S0(n345) );
  HS65_GSS_XNOR2X3 U280 ( .A(n349), .B(n348), .Z(n870) );
  HS65_GS_IVX2 U281 ( .A(n870), .Z(n347) );
  HS65_GS_AOI12X2 U282 ( .A(n344), .B(n345), .C(n347), .Z(n869) );
  HS65_GS_NAND2X2 U283 ( .A(n345), .B(n344), .Z(n343) );
  HS65_GS_IVX2 U284 ( .A(n343), .Z(n346) );
  HS65_GS_AND2X4 U285 ( .A(\mul_b0/fa1_s0_r[28] ), .B(\mul_b0/fa1_s1_r[28] ), 
        .Z(n246) );
  HS65_GSS_XOR2X3 U286 ( .A(\mul_b0/fa1_s0_r[29] ), .B(\mul_b0/fa1_s1_r[29] ), 
        .Z(n245) );
  HS65_GS_FA1X4 U287 ( .A0(\mul_b0/fa1_s2_r[30] ), .B0(n244), .CI(n243), .CO(
        n344), .S0(n880) );
  HS65_GS_AND2X4 U288 ( .A(\mul_b0/fa1_s0_r[27] ), .B(\mul_b0/fa1_s1_r[27] ), 
        .Z(n248) );
  HS65_GSS_XOR2X3 U289 ( .A(\mul_b0/fa1_s0_r[28] ), .B(\mul_b0/fa1_s1_r[28] ), 
        .Z(n247) );
  HS65_GS_FA1X4 U290 ( .A0(\mul_b0/fa1_s2_r[29] ), .B0(n246), .CI(n245), .CO(
        n881), .S0(n877) );
  HS65_GS_AND2X4 U291 ( .A(\mul_b0/fa1_s0_r[26] ), .B(\mul_b0/fa1_s1_r[26] ), 
        .Z(n336) );
  HS65_GSS_XOR2X3 U292 ( .A(\mul_b0/fa1_s0_r[27] ), .B(\mul_b0/fa1_s1_r[27] ), 
        .Z(n335) );
  HS65_GS_FA1X4 U293 ( .A0(\mul_b0/fa1_s2_r[28] ), .B0(n248), .CI(n247), .CO(
        n878), .S0(n1051) );
  HS65_GSS_XOR2X3 U294 ( .A(\mul_b0/fa1_s0_r[25] ), .B(\mul_b0/fa1_s1_r[25] ), 
        .Z(n250) );
  HS65_GS_AND2X4 U295 ( .A(\mul_b0/fa1_s0_r[24] ), .B(\mul_b0/fa1_s1_r[24] ), 
        .Z(n249) );
  HS65_GS_AND2X4 U296 ( .A(\mul_b0/fa1_s1_r[25] ), .B(\mul_b0/fa1_s0_r[25] ), 
        .Z(n338) );
  HS65_GSS_XOR2X3 U297 ( .A(\mul_b0/fa1_s0_r[26] ), .B(\mul_b0/fa1_s1_r[26] ), 
        .Z(n337) );
  HS65_GS_AND2X4 U298 ( .A(\mul_b0/fa1_s0_r[23] ), .B(\mul_b0/fa1_s1_r[23] ), 
        .Z(n252) );
  HS65_GSS_XOR2X3 U299 ( .A(\mul_b0/fa1_s0_r[24] ), .B(\mul_b0/fa1_s1_r[24] ), 
        .Z(n251) );
  HS65_GS_FA1X4 U300 ( .A0(\mul_b0/fa1_s2_r[25] ), .B0(n250), .CI(n249), .CO(
        n334), .S0(n330) );
  HS65_GS_AND2X4 U301 ( .A(\mul_b0/fa1_s0_r[22] ), .B(\mul_b0/fa1_s1_r[22] ), 
        .Z(n254) );
  HS65_GSS_XOR2X3 U302 ( .A(\mul_b0/fa1_s0_r[23] ), .B(\mul_b0/fa1_s1_r[23] ), 
        .Z(n253) );
  HS65_GS_FA1X4 U303 ( .A0(\mul_b0/fa1_s2_r[24] ), .B0(n252), .CI(n251), .CO(
        n331), .S0(n327) );
  HS65_GSS_XOR2X3 U304 ( .A(\mul_b0/fa1_s0_r[22] ), .B(\mul_b0/fa1_s1_r[22] ), 
        .Z(n255) );
  HS65_GS_FA1X4 U305 ( .A0(\mul_b0/fa1_s2_r[23] ), .B0(n254), .CI(n253), .CO(
        n328), .S0(n324) );
  HS65_GS_FA1X4 U306 ( .A0(\mul_b0/fa1_s0_r[21] ), .B0(\mul_b0/fa1_s1_r[21] ), 
        .CI(\mul_b0/fa1_c0_r[20] ), .CO(n256), .S0(n258) );
  HS65_GS_FA1X4 U307 ( .A0(\mul_b0/fa1_s2_r[22] ), .B0(n256), .CI(n255), .CO(
        n325), .S0(n321) );
  HS65_GS_FA1X4 U308 ( .A0(\mul_b0/fa1_s0_r[20] ), .B0(\mul_b0/fa1_s1_r[20] ), 
        .CI(\mul_b0/fa1_c0_r[19] ), .CO(n257), .S0(n259) );
  HS65_GS_FA1X4 U309 ( .A0(\mul_b0/fa1_s2_r[21] ), .B0(n258), .CI(n257), .CO(
        n322), .S0(n318) );
  HS65_GS_FA1X4 U310 ( .A0(\mul_b0/fa1_s0_r[19] ), .B0(\mul_b0/fa1_s1_r[19] ), 
        .CI(\mul_b0/fa1_c0_r[18] ), .CO(n260), .S0(n261) );
  HS65_GS_FA1X4 U311 ( .A0(\mul_b0/fa1_s2_r[20] ), .B0(n260), .CI(n259), .CO(
        n319), .S0(n315) );
  HS65_GS_FA1X4 U312 ( .A0(\mul_b0/fa1_s0_r[18] ), .B0(\mul_b0/fa1_s1_r[18] ), 
        .CI(\mul_b0/fa1_c0_r[17] ), .CO(n262), .S0(n263) );
  HS65_GS_FA1X4 U313 ( .A0(\mul_b0/fa1_s2_r[19] ), .B0(n262), .CI(n261), .CO(
        n316), .S0(n312) );
  HS65_GS_FA1X4 U314 ( .A0(\mul_b0/fa1_s0_r[17] ), .B0(\mul_b0/fa1_s1_r[17] ), 
        .CI(\mul_b0/fa1_c0_r[16] ), .CO(n264), .S0(n265) );
  HS65_GS_FA1X4 U315 ( .A0(\mul_b0/fa1_s2_r[18] ), .B0(n264), .CI(n263), .CO(
        n313), .S0(n309) );
  HS65_GS_FA1X4 U316 ( .A0(\mul_b0/fa1_s0_r[16] ), .B0(\mul_b0/fa1_s1_r[16] ), 
        .CI(\mul_b0/fa1_c0_r[15] ), .CO(n266), .S0(n267) );
  HS65_GS_FA1X4 U317 ( .A0(\mul_b0/fa1_s2_r[17] ), .B0(n266), .CI(n265), .CO(
        n310), .S0(n306) );
  HS65_GS_FA1X4 U318 ( .A0(\mul_b0/fa1_s0_r[15] ), .B0(\mul_b0/fa1_s1_r[15] ), 
        .CI(\mul_b0/fa1_c0_r[14] ), .CO(n268), .S0(n271) );
  HS65_GS_FA1X4 U319 ( .A0(\mul_b0/fa1_s2_r[16] ), .B0(n268), .CI(n267), .CO(
        n307), .S0(n303) );
  HS65_GS_NOR2X2 U320 ( .A(n304), .B(n303), .Z(n269) );
  HS65_GS_AOI12X2 U321 ( .A(n303), .B(n304), .C(n269), .Z(n930) );
  HS65_GS_FA1X4 U322 ( .A0(\mul_b0/fa1_s0_r[14] ), .B0(\mul_b0/fa1_s1_r[14] ), 
        .CI(\mul_b0/fa1_c0_r[13] ), .CO(n270), .S0(n273) );
  HS65_GS_FA1X4 U323 ( .A0(\mul_b0/fa1_s2_r[15] ), .B0(n271), .CI(n270), .CO(
        n304), .S0(n300) );
  HS65_GS_FA1X4 U324 ( .A0(\mul_b0/fa1_s0_r[13] ), .B0(\mul_b0/fa1_s1_r[13] ), 
        .CI(\mul_b0/fa1_c0_r[12] ), .CO(n272), .S0(n274) );
  HS65_GS_FA1X4 U325 ( .A0(\mul_b0/fa1_s2_r[14] ), .B0(n273), .CI(n272), .CO(
        n301), .S0(n297) );
  HS65_GS_FA1X4 U326 ( .A0(\mul_b0/fa1_s0_r[12] ), .B0(\mul_b0/fa1_s1_r[12] ), 
        .CI(\mul_b0/fa1_c0_r[11] ), .CO(n275), .S0(n287) );
  HS65_GS_FA1X4 U327 ( .A0(\mul_b0/fa1_s2_r[13] ), .B0(n275), .CI(n274), .CO(
        n298), .S0(n294) );
  HS65_GS_FA1X4 U328 ( .A0(\mul_b0/fa1_s0_r[11] ), .B0(\mul_b0/fa1_s1_r[11] ), 
        .CI(\mul_b0/fa1_c0_r[10] ), .CO(n288), .S0(n292) );
  HS65_GS_NOR2X2 U329 ( .A(n291), .B(n292), .Z(n286) );
  HS65_GS_FA1X4 U330 ( .A0(\mul_b0/fa1_s0_r[10] ), .B0(\mul_b0/fa1_s1_r[10] ), 
        .CI(\mul_b0/fa1_c0_r[9] ), .CO(n291), .S0(n284) );
  HS65_GS_FA1X4 U331 ( .A0(\mul_b0/fa1_s0_r[9] ), .B0(\mul_b0/fa1_s1_r[9] ), 
        .CI(\mul_b0/fa1_c0_r[8] ), .CO(n283), .S0(n281) );
  HS65_GS_FA1X4 U332 ( .A0(\mul_b0/fa1_s0_r[8] ), .B0(\mul_b0/fa1_s1_r[8] ), 
        .CI(\mul_b0/fa1_c0_r[7] ), .CO(n280), .S0(n278) );
  HS65_GS_AND2X4 U333 ( .A(\mul_b0/fa1_s0_r[6] ), .B(\mul_b0/fa1_c0_r[5] ), 
        .Z(n276) );
  HS65_GS_PAOI2X1 U334 ( .A(\mul_b0/fa1_c0_r[6] ), .B(n276), .P(
        \mul_b0/fa1_s0_r[7] ), .Z(n277) );
  HS65_GS_NOR2AX3 U335 ( .A(n278), .B(n277), .Z(n279) );
  HS65_GS_PAO2X4 U336 ( .A(n281), .B(n280), .P(n279), .Z(n282) );
  HS65_GS_PAOI2X1 U337 ( .A(n284), .B(n283), .P(n282), .Z(n285) );
  HS65_GS_NOR2X2 U338 ( .A(n286), .B(n285), .Z(n290) );
  HS65_GS_FA1X4 U339 ( .A0(\mul_b0/fa1_s2_r[12] ), .B0(n288), .CI(n287), .CO(
        n295), .S0(n289) );
  HS65_GS_CB4I1X4 U340 ( .A(n292), .B(n291), .C(n290), .D(n289), .Z(n293) );
  HS65_GS_PAOI2X1 U341 ( .A(n295), .B(n294), .P(n293), .Z(n937) );
  HS65_GS_NAND2X2 U342 ( .A(n297), .B(n298), .Z(n296) );
  HS65_GS_OAI21X2 U343 ( .A(n297), .B(n298), .C(n296), .Z(n936) );
  HS65_GS_NOR2X2 U344 ( .A(n937), .B(n936), .Z(n935) );
  HS65_GS_AOI12X2 U345 ( .A(n298), .B(n297), .C(n935), .Z(n933) );
  HS65_GS_NAND2X2 U346 ( .A(n300), .B(n301), .Z(n299) );
  HS65_GS_OAI21X2 U347 ( .A(n300), .B(n301), .C(n299), .Z(n932) );
  HS65_GS_NOR2X2 U348 ( .A(n933), .B(n932), .Z(n931) );
  HS65_GS_AOI12X2 U349 ( .A(n301), .B(n300), .C(n931), .Z(n929) );
  HS65_GS_NAND2X2 U350 ( .A(n930), .B(n929), .Z(n302) );
  HS65_GS_OAI21X2 U351 ( .A(n304), .B(n303), .C(n302), .Z(n926) );
  HS65_GS_NAND2X2 U352 ( .A(n306), .B(n307), .Z(n305) );
  HS65_GS_OAI21X2 U353 ( .A(n306), .B(n307), .C(n305), .Z(n925) );
  HS65_GS_NOR2X2 U354 ( .A(n926), .B(n925), .Z(n924) );
  HS65_GS_AOI12X2 U355 ( .A(n307), .B(n306), .C(n924), .Z(n922) );
  HS65_GS_NAND2X2 U356 ( .A(n309), .B(n310), .Z(n308) );
  HS65_GS_OAI21X2 U357 ( .A(n309), .B(n310), .C(n308), .Z(n921) );
  HS65_GS_NOR2X2 U358 ( .A(n922), .B(n921), .Z(n920) );
  HS65_GS_AOI12X2 U359 ( .A(n310), .B(n309), .C(n920), .Z(n918) );
  HS65_GS_NAND2X2 U360 ( .A(n312), .B(n313), .Z(n311) );
  HS65_GS_OAI21X2 U361 ( .A(n312), .B(n313), .C(n311), .Z(n917) );
  HS65_GS_NOR2X2 U362 ( .A(n918), .B(n917), .Z(n916) );
  HS65_GS_AOI12X2 U363 ( .A(n313), .B(n312), .C(n916), .Z(n914) );
  HS65_GS_NAND2X2 U364 ( .A(n315), .B(n316), .Z(n314) );
  HS65_GS_OAI21X2 U365 ( .A(n315), .B(n316), .C(n314), .Z(n913) );
  HS65_GS_NOR2X2 U366 ( .A(n914), .B(n913), .Z(n912) );
  HS65_GS_AOI12X2 U367 ( .A(n316), .B(n315), .C(n912), .Z(n910) );
  HS65_GS_NAND2X2 U368 ( .A(n318), .B(n319), .Z(n317) );
  HS65_GS_OAI21X2 U369 ( .A(n318), .B(n319), .C(n317), .Z(n909) );
  HS65_GS_NOR2X2 U370 ( .A(n910), .B(n909), .Z(n908) );
  HS65_GS_AOI12X2 U371 ( .A(n319), .B(n318), .C(n908), .Z(n906) );
  HS65_GS_NAND2X2 U372 ( .A(n321), .B(n322), .Z(n320) );
  HS65_GS_OAI21X2 U373 ( .A(n321), .B(n322), .C(n320), .Z(n905) );
  HS65_GS_NOR2X2 U374 ( .A(n906), .B(n905), .Z(n904) );
  HS65_GS_AOI12X2 U375 ( .A(n322), .B(n321), .C(n904), .Z(n902) );
  HS65_GS_NAND2X2 U376 ( .A(n324), .B(n325), .Z(n323) );
  HS65_GS_OAI21X2 U377 ( .A(n324), .B(n325), .C(n323), .Z(n901) );
  HS65_GS_NOR2X2 U378 ( .A(n902), .B(n901), .Z(n900) );
  HS65_GS_AOI12X2 U379 ( .A(n325), .B(n324), .C(n900), .Z(n898) );
  HS65_GS_NAND2X2 U380 ( .A(n327), .B(n328), .Z(n326) );
  HS65_GS_OAI21X2 U381 ( .A(n327), .B(n328), .C(n326), .Z(n897) );
  HS65_GS_NOR2X2 U382 ( .A(n898), .B(n897), .Z(n896) );
  HS65_GS_AOI12X2 U383 ( .A(n328), .B(n327), .C(n896), .Z(n894) );
  HS65_GS_NAND2X2 U384 ( .A(n330), .B(n331), .Z(n329) );
  HS65_GS_OAI21X2 U385 ( .A(n330), .B(n331), .C(n329), .Z(n893) );
  HS65_GS_NOR2X2 U386 ( .A(n894), .B(n893), .Z(n892) );
  HS65_GS_AOI12X2 U387 ( .A(n331), .B(n330), .C(n892), .Z(n890) );
  HS65_GS_NAND2X2 U388 ( .A(n333), .B(n334), .Z(n332) );
  HS65_GS_OAI21X2 U389 ( .A(n333), .B(n334), .C(n332), .Z(n889) );
  HS65_GS_NOR2X2 U390 ( .A(n890), .B(n889), .Z(n888) );
  HS65_GS_AOI12X2 U391 ( .A(n334), .B(n333), .C(n888), .Z(n1058) );
  HS65_GS_FA1X4 U392 ( .A0(\mul_b0/fa1_s2_r[27] ), .B0(n336), .CI(n335), .CO(
        n1052), .S0(n340) );
  HS65_GS_FA1X4 U393 ( .A0(\mul_b0/fa1_s2_r[26] ), .B0(n338), .CI(n337), .CO(
        n339), .S0(n333) );
  HS65_GS_NAND2X2 U394 ( .A(n340), .B(n339), .Z(n341) );
  HS65_GS_OAI21X2 U395 ( .A(n340), .B(n339), .C(n341), .Z(n1059) );
  HS65_GS_OAI21X2 U396 ( .A(n1058), .B(n1059), .C(n341), .Z(n1050) );
  HS65_GS_IVX2 U397 ( .A(n342), .Z(n875) );
  HS65_GS_OAI21X2 U398 ( .A(n345), .B(n344), .C(n343), .Z(n874) );
  HS65_GS_NOR2X2 U399 ( .A(n875), .B(n874), .Z(n873) );
  HS65_GS_AOI12X2 U400 ( .A(n347), .B(n346), .C(n873), .Z(n872) );
  HS65_GS_NAND2X2 U401 ( .A(n349), .B(n348), .Z(n350) );
  HS65_GS_OAI21X2 U402 ( .A(n869), .B(n872), .C(n350), .Z(n351) );
  HS65_GSS_XOR3X2 U403 ( .A(n353), .B(n352), .C(n351), .Z(n354) );
  HS65_GSS_XOR2X3 U404 ( .A(\mul_b0/fa1_s2_r[33] ), .B(n354), .Z(n355) );
  HS65_GSS_XOR3X2 U405 ( .A(\mul_b0/fa1_s0_r[33] ), .B(\mul_b0/fa1_s1_r[33] ), 
        .C(n355), .Z(\mul_b0/result_sat[15] ) );
  HS65_GS_AND2X4 U406 ( .A(\mul_b1/fa1_c2_r[28] ), .B(\mul_b1/fa1_s2_r[29] ), 
        .Z(n515) );
  HS65_GSS_XOR2X3 U407 ( .A(\mul_b1/fa1_s2_r[29] ), .B(\mul_b1/fa1_c2_r[28] ), 
        .Z(n506) );
  HS65_GSS_XOR2X3 U408 ( .A(\mul_b1/fa1_s1_r[29] ), .B(\mul_b1/fa1_s0_r[29] ), 
        .Z(n505) );
  HS65_GS_AND2X4 U409 ( .A(\mul_b1/fa1_s1_r[28] ), .B(\mul_b1/fa1_s0_r[28] ), 
        .Z(n504) );
  HS65_GS_AND2X4 U410 ( .A(\mul_b1/fa1_s1_r[29] ), .B(\mul_b1/fa1_s0_r[29] ), 
        .Z(n517) );
  HS65_GSS_XOR2X3 U411 ( .A(\mul_b1/fa1_s1_r[30] ), .B(\mul_b1/fa1_s0_r[30] ), 
        .Z(n516) );
  HS65_GS_AND2X4 U412 ( .A(\mul_b1/fa1_c2_r[26] ), .B(\mul_b1/fa1_s2_r[27] ), 
        .Z(n503) );
  HS65_GSS_XOR2X3 U413 ( .A(\mul_b1/fa1_s2_r[27] ), .B(\mul_b1/fa1_c2_r[26] ), 
        .Z(n358) );
  HS65_GSS_XOR2X3 U414 ( .A(\mul_b1/fa1_s1_r[27] ), .B(\mul_b1/fa1_s0_r[27] ), 
        .Z(n357) );
  HS65_GS_AND2X4 U415 ( .A(\mul_b1/fa1_s0_r[26] ), .B(\mul_b1/fa1_s1_r[26] ), 
        .Z(n356) );
  HS65_GS_AND2X4 U416 ( .A(\mul_b1/fa1_s1_r[27] ), .B(\mul_b1/fa1_s0_r[27] ), 
        .Z(n509) );
  HS65_GSS_XOR2X3 U417 ( .A(\mul_b1/fa1_s2_r[28] ), .B(\mul_b1/fa1_c2_r[27] ), 
        .Z(n508) );
  HS65_GSS_XOR2X3 U418 ( .A(\mul_b1/fa1_s1_r[28] ), .B(\mul_b1/fa1_s0_r[28] ), 
        .Z(n507) );
  HS65_GS_AND2X4 U419 ( .A(\mul_b1/fa1_c2_r[25] ), .B(\mul_b1/fa1_s2_r[26] ), 
        .Z(n500) );
  HS65_GSS_XOR2X3 U420 ( .A(\mul_b1/fa1_s2_r[26] ), .B(\mul_b1/fa1_c2_r[25] ), 
        .Z(n491) );
  HS65_GSS_XOR2X3 U421 ( .A(\mul_b1/fa1_s0_r[26] ), .B(\mul_b1/fa1_s1_r[26] ), 
        .Z(n490) );
  HS65_GS_AND2X4 U422 ( .A(\mul_b1/fa1_s0_r[25] ), .B(\mul_b1/fa1_s1_r[25] ), 
        .Z(n489) );
  HS65_GS_FA1X4 U423 ( .A0(n358), .B0(n357), .CI(n356), .CO(n502), .S0(n498)
         );
  HS65_GS_AND2X4 U424 ( .A(\mul_b1/fa1_c2_r[23] ), .B(\mul_b1/fa1_s2_r[24] ), 
        .Z(n488) );
  HS65_GSS_XOR2X3 U425 ( .A(\mul_b1/fa1_s2_r[24] ), .B(\mul_b1/fa1_c2_r[23] ), 
        .Z(n361) );
  HS65_GSS_XOR2X3 U426 ( .A(\mul_b1/fa1_s1_r[24] ), .B(\mul_b1/fa1_s0_r[24] ), 
        .Z(n360) );
  HS65_GS_AND2X4 U427 ( .A(\mul_b1/fa1_s0_r[23] ), .B(\mul_b1/fa1_s1_r[23] ), 
        .Z(n359) );
  HS65_GS_AND2X4 U428 ( .A(\mul_b1/fa1_s1_r[24] ), .B(\mul_b1/fa1_s0_r[24] ), 
        .Z(n494) );
  HS65_GSS_XOR2X3 U429 ( .A(\mul_b1/fa1_s2_r[25] ), .B(\mul_b1/fa1_c2_r[24] ), 
        .Z(n493) );
  HS65_GSS_XOR2X3 U430 ( .A(\mul_b1/fa1_s0_r[25] ), .B(\mul_b1/fa1_s1_r[25] ), 
        .Z(n492) );
  HS65_GS_FA1X4 U431 ( .A0(\mul_b1/fa1_c1_r[22] ), .B0(\mul_b1/fa1_c2_r[22] ), 
        .CI(\mul_b1/fa1_s2_r[23] ), .CO(n485), .S0(n364) );
  HS65_GSS_XOR2X3 U432 ( .A(\mul_b1/fa1_s0_r[23] ), .B(\mul_b1/fa1_s1_r[23] ), 
        .Z(n363) );
  HS65_GS_AND2X4 U433 ( .A(\mul_b1/fa1_s0_r[22] ), .B(\mul_b1/fa1_s1_r[22] ), 
        .Z(n362) );
  HS65_GS_FA1X4 U434 ( .A0(n361), .B0(n360), .CI(n359), .CO(n487), .S0(n483)
         );
  HS65_GS_FA1X4 U435 ( .A0(\mul_b1/fa1_c1_r[21] ), .B0(\mul_b1/fa1_c2_r[21] ), 
        .CI(\mul_b1/fa1_s2_r[22] ), .CO(n367), .S0(n479) );
  HS65_GSS_XOR2X3 U436 ( .A(\mul_b1/fa1_s0_r[22] ), .B(\mul_b1/fa1_s1_r[22] ), 
        .Z(n478) );
  HS65_GS_AND2X4 U437 ( .A(\mul_b1/fa1_s1_r[21] ), .B(\mul_b1/fa1_s0_r[21] ), 
        .Z(n477) );
  HS65_GS_FA1X4 U438 ( .A0(n364), .B0(n363), .CI(n362), .CO(n484), .S0(n365)
         );
  HS65_GS_FA1X4 U439 ( .A0(n367), .B0(n366), .CI(n365), .CO(n1118), .S0(n1125)
         );
  HS65_GS_AND2X4 U440 ( .A(\mul_b1/fa1_c1_r[13] ), .B(\mul_b1/fa1_s2_r[14] ), 
        .Z(n419) );
  HS65_GSS_XOR2X3 U441 ( .A(\mul_b1/fa1_s1_r[15] ), .B(\mul_b1/fa1_s0_r[15] ), 
        .Z(n421) );
  HS65_GS_AND2X4 U442 ( .A(\mul_b1/fa1_s1_r[14] ), .B(\mul_b1/fa1_s0_r[14] ), 
        .Z(n420) );
  HS65_GSS_XOR2X3 U443 ( .A(\mul_b1/fa1_s1_r[14] ), .B(\mul_b1/fa1_s0_r[14] ), 
        .Z(n370) );
  HS65_GSS_XOR2X3 U444 ( .A(\mul_b1/fa1_c1_r[13] ), .B(\mul_b1/fa1_s2_r[14] ), 
        .Z(n369) );
  HS65_GS_AND2X4 U445 ( .A(\mul_b1/fa1_s1_r[13] ), .B(\mul_b1/fa1_s0_r[13] ), 
        .Z(n368) );
  HS65_GS_IVX2 U446 ( .A(n414), .Z(n416) );
  HS65_GS_AND2X4 U447 ( .A(\mul_b1/fa1_s2_r[13] ), .B(\mul_b1/fa1_c1_r[12] ), 
        .Z(n413) );
  HS65_GS_FA1X4 U448 ( .A0(n370), .B0(n369), .CI(n368), .CO(n417), .S0(n412)
         );
  HS65_GS_AND2X4 U449 ( .A(\mul_b1/fa1_s0_r[12] ), .B(\mul_b1/fa1_s1_r[12] ), 
        .Z(n401) );
  HS65_GSS_XOR2X3 U450 ( .A(\mul_b1/fa1_s2_r[13] ), .B(\mul_b1/fa1_c1_r[12] ), 
        .Z(n400) );
  HS65_GSS_XOR2X3 U451 ( .A(\mul_b1/fa1_s1_r[13] ), .B(\mul_b1/fa1_s0_r[13] ), 
        .Z(n399) );
  HS65_GSS_XOR2X3 U452 ( .A(\mul_b1/fa1_s0_r[12] ), .B(\mul_b1/fa1_s1_r[12] ), 
        .Z(n403) );
  HS65_GS_AND2X4 U453 ( .A(\mul_b1/fa1_s0_r[11] ), .B(\mul_b1/fa1_s1_r[11] ), 
        .Z(n402) );
  HS65_GSS_XOR2X3 U454 ( .A(\mul_b1/fa1_s0_r[11] ), .B(\mul_b1/fa1_s1_r[11] ), 
        .Z(n372) );
  HS65_GS_AND2X4 U455 ( .A(\mul_b1/fa1_s0_r[10] ), .B(\mul_b1/fa1_s1_r[10] ), 
        .Z(n371) );
  HS65_GSS_XOR2X3 U456 ( .A(n397), .B(n398), .Z(n396) );
  HS65_GSS_XOR2X3 U457 ( .A(\mul_b1/fa1_s0_r[10] ), .B(\mul_b1/fa1_s1_r[10] ), 
        .Z(n374) );
  HS65_GS_AND2X4 U458 ( .A(\mul_b1/fa1_s0_r[9] ), .B(\mul_b1/fa1_s1_r[9] ), 
        .Z(n373) );
  HS65_GS_FA1X4 U459 ( .A0(\mul_b1/fa1_c1_r[10] ), .B0(n372), .CI(n371), .CO(
        n398), .S0(n389) );
  HS65_GS_AND2X4 U460 ( .A(n388), .B(n389), .Z(n395) );
  HS65_GS_FA1X4 U461 ( .A0(\mul_b1/fa1_c1_r[9] ), .B0(n374), .CI(n373), .CO(
        n388), .S0(n386) );
  HS65_GS_IVX2 U462 ( .A(n386), .Z(n393) );
  HS65_GS_NAND2X2 U463 ( .A(\mul_b1/fa1_s1_r[7] ), .B(\mul_b1/fa1_s0_r[7] ), 
        .Z(n375) );
  HS65_GSS_XNOR2X3 U464 ( .A(\mul_b1/fa1_s0_r[8] ), .B(\mul_b1/fa1_s1_r[8] ), 
        .Z(n378) );
  HS65_GS_NOR2X2 U465 ( .A(n375), .B(n378), .Z(n383) );
  HS65_GSS_XOR2X3 U466 ( .A(\mul_b1/fa1_s0_r[9] ), .B(\mul_b1/fa1_s1_r[9] ), 
        .Z(n385) );
  HS65_GS_AND2X4 U467 ( .A(\mul_b1/fa1_s0_r[8] ), .B(\mul_b1/fa1_s1_r[8] ), 
        .Z(n384) );
  HS65_GS_NAND2X2 U468 ( .A(\mul_b1/fa1_s1_r[6] ), .B(\mul_b1/fa1_s0_r[6] ), 
        .Z(n377) );
  HS65_GSS_XNOR2X3 U469 ( .A(\mul_b1/fa1_s1_r[7] ), .B(\mul_b1/fa1_s0_r[7] ), 
        .Z(n376) );
  HS65_GS_NOR2X2 U470 ( .A(n377), .B(n376), .Z(n380) );
  HS65_GS_IVX2 U471 ( .A(n378), .Z(n379) );
  HS65_GS_AND2X4 U472 ( .A(n380), .B(n379), .Z(n381) );
  HS65_GS_PAOI2X1 U473 ( .A(n383), .B(n382), .P(n381), .Z(n392) );
  HS65_GS_FA1X4 U474 ( .A0(\mul_b1/fa1_c1_r[8] ), .B0(n385), .CI(n384), .CO(
        n387), .S0(n382) );
  HS65_GS_NAND2X2 U475 ( .A(n387), .B(n386), .Z(n391) );
  HS65_GSS_XNOR2X3 U476 ( .A(n389), .B(n388), .Z(n390) );
  HS65_GS_CBI4I6X2 U477 ( .A(n393), .B(n392), .C(n391), .D(n390), .Z(n394) );
  HS65_GS_PAO2X4 U478 ( .A(n396), .B(n395), .P(n394), .Z(n406) );
  HS65_GS_AND2X4 U479 ( .A(n398), .B(n397), .Z(n405) );
  HS65_GS_FA1X4 U480 ( .A0(n401), .B0(n400), .CI(n399), .CO(n411), .S0(n407)
         );
  HS65_GS_FA1X4 U481 ( .A0(\mul_b1/fa1_c1_r[11] ), .B0(n403), .CI(n402), .CO(
        n408), .S0(n397) );
  HS65_GSS_XOR2X3 U482 ( .A(n407), .B(n408), .Z(n404) );
  HS65_GS_PAOI2X1 U483 ( .A(n406), .B(n405), .P(n404), .Z(n410) );
  HS65_GS_AND2X4 U484 ( .A(n408), .B(n407), .Z(n409) );
  HS65_GS_NOR2AX3 U485 ( .A(n410), .B(n409), .Z(n1748) );
  HS65_GS_FA1X4 U486 ( .A0(n413), .B0(n412), .CI(n411), .CO(n1754), .S0(n1749)
         );
  HS65_GS_NOR2X2 U487 ( .A(n1749), .B(n1748), .Z(n1747) );
  HS65_GS_NOR2X2 U488 ( .A(n1748), .B(n1747), .Z(n415) );
  HS65_GSS_XNOR2X3 U489 ( .A(n415), .B(n414), .Z(n1753) );
  HS65_GS_NOR2X2 U490 ( .A(n1754), .B(n1753), .Z(n1752) );
  HS65_GS_NOR2X2 U491 ( .A(n416), .B(n1752), .Z(n424) );
  HS65_GS_FA1X4 U492 ( .A0(n419), .B0(n418), .CI(n417), .CO(n423), .S0(n414)
         );
  HS65_GS_NOR2X2 U493 ( .A(n424), .B(n423), .Z(n425) );
  HS65_GS_FA1X4 U494 ( .A0(\mul_b1/fa1_c1_r[14] ), .B0(\mul_b1/fa1_c2_r[14] ), 
        .CI(\mul_b1/fa1_s2_r[15] ), .CO(n428), .S0(n422) );
  HS65_GS_FA1X4 U495 ( .A0(n422), .B0(n421), .CI(n420), .CO(n427), .S0(n418)
         );
  HS65_GSS_XOR2X3 U496 ( .A(\mul_b1/fa1_s1_r[16] ), .B(\mul_b1/fa1_s0_r[16] ), 
        .Z(n430) );
  HS65_GS_AND2X4 U497 ( .A(\mul_b1/fa1_s1_r[15] ), .B(\mul_b1/fa1_s0_r[15] ), 
        .Z(n429) );
  HS65_GSS_XNOR2X3 U498 ( .A(n424), .B(n423), .Z(n1757) );
  HS65_GS_NOR2X2 U499 ( .A(n1758), .B(n1757), .Z(n1756) );
  HS65_GS_NOR2X2 U500 ( .A(n425), .B(n1756), .Z(n433) );
  HS65_GS_FA1X4 U501 ( .A0(n428), .B0(n427), .CI(n426), .CO(n432), .S0(n1758)
         );
  HS65_GS_NOR2X2 U502 ( .A(n433), .B(n432), .Z(n434) );
  HS65_GS_FA1X4 U503 ( .A0(\mul_b1/fa1_c1_r[15] ), .B0(\mul_b1/fa1_c2_r[15] ), 
        .CI(\mul_b1/fa1_s2_r[16] ), .CO(n437), .S0(n431) );
  HS65_GS_FA1X4 U504 ( .A0(n431), .B0(n430), .CI(n429), .CO(n436), .S0(n426)
         );
  HS65_GSS_XOR2X3 U505 ( .A(\mul_b1/fa1_s1_r[17] ), .B(\mul_b1/fa1_s0_r[17] ), 
        .Z(n439) );
  HS65_GS_AND2X4 U506 ( .A(\mul_b1/fa1_s1_r[16] ), .B(\mul_b1/fa1_s0_r[16] ), 
        .Z(n438) );
  HS65_GSS_XNOR2X3 U507 ( .A(n433), .B(n432), .Z(n1761) );
  HS65_GS_NOR2X2 U508 ( .A(n1762), .B(n1761), .Z(n1760) );
  HS65_GS_NOR2X2 U509 ( .A(n434), .B(n1760), .Z(n441) );
  HS65_GS_FA1X4 U510 ( .A0(n437), .B0(n436), .CI(n435), .CO(n442), .S0(n1762)
         );
  HS65_GS_NOR2X2 U511 ( .A(n441), .B(n442), .Z(n443) );
  HS65_GS_FA1X4 U512 ( .A0(\mul_b1/fa1_c1_r[16] ), .B0(\mul_b1/fa1_c2_r[16] ), 
        .CI(\mul_b1/fa1_s2_r[17] ), .CO(n446), .S0(n440) );
  HS65_GS_FA1X4 U513 ( .A0(n440), .B0(n439), .CI(n438), .CO(n445), .S0(n435)
         );
  HS65_GSS_XOR2X3 U514 ( .A(\mul_b1/fa1_s1_r[18] ), .B(\mul_b1/fa1_s0_r[18] ), 
        .Z(n448) );
  HS65_GS_AND2X4 U515 ( .A(\mul_b1/fa1_s1_r[17] ), .B(\mul_b1/fa1_s0_r[17] ), 
        .Z(n447) );
  HS65_GSS_XNOR2X3 U516 ( .A(n442), .B(n441), .Z(n1765) );
  HS65_GS_NOR2X2 U517 ( .A(n1766), .B(n1765), .Z(n1764) );
  HS65_GS_NOR2X2 U518 ( .A(n443), .B(n1764), .Z(n450) );
  HS65_GS_FA1X4 U519 ( .A0(n446), .B0(n445), .CI(n444), .CO(n451), .S0(n1766)
         );
  HS65_GS_NOR2X2 U520 ( .A(n450), .B(n451), .Z(n452) );
  HS65_GS_FA1X4 U521 ( .A0(\mul_b1/fa1_c1_r[17] ), .B0(\mul_b1/fa1_c2_r[17] ), 
        .CI(\mul_b1/fa1_s2_r[18] ), .CO(n455), .S0(n449) );
  HS65_GS_FA1X4 U522 ( .A0(n449), .B0(n448), .CI(n447), .CO(n454), .S0(n444)
         );
  HS65_GSS_XOR2X3 U523 ( .A(\mul_b1/fa1_s1_r[19] ), .B(\mul_b1/fa1_s0_r[19] ), 
        .Z(n457) );
  HS65_GS_AND2X4 U524 ( .A(\mul_b1/fa1_s1_r[18] ), .B(\mul_b1/fa1_s0_r[18] ), 
        .Z(n456) );
  HS65_GSS_XNOR2X3 U525 ( .A(n451), .B(n450), .Z(n1769) );
  HS65_GS_NOR2X2 U526 ( .A(n1770), .B(n1769), .Z(n1768) );
  HS65_GS_NOR2X2 U527 ( .A(n452), .B(n1768), .Z(n459) );
  HS65_GS_FA1X4 U528 ( .A0(n455), .B0(n454), .CI(n453), .CO(n460), .S0(n1770)
         );
  HS65_GS_NOR2X2 U529 ( .A(n459), .B(n460), .Z(n461) );
  HS65_GS_FA1X4 U530 ( .A0(\mul_b1/fa1_c1_r[18] ), .B0(\mul_b1/fa1_c2_r[18] ), 
        .CI(\mul_b1/fa1_s2_r[19] ), .CO(n464), .S0(n458) );
  HS65_GS_FA1X4 U531 ( .A0(n458), .B0(n457), .CI(n456), .CO(n463), .S0(n453)
         );
  HS65_GSS_XOR2X3 U532 ( .A(\mul_b1/fa1_s1_r[20] ), .B(\mul_b1/fa1_s0_r[20] ), 
        .Z(n467) );
  HS65_GS_AND2X4 U533 ( .A(\mul_b1/fa1_s1_r[19] ), .B(\mul_b1/fa1_s0_r[19] ), 
        .Z(n465) );
  HS65_GSS_XNOR2X3 U534 ( .A(n460), .B(n459), .Z(n1773) );
  HS65_GS_NOR2X2 U535 ( .A(n1774), .B(n1773), .Z(n1772) );
  HS65_GS_NOR2X2 U536 ( .A(n461), .B(n1772), .Z(n468) );
  HS65_GS_FA1X4 U537 ( .A0(n464), .B0(n463), .CI(n462), .CO(n469), .S0(n1774)
         );
  HS65_GS_NOR2X2 U538 ( .A(n468), .B(n469), .Z(n470) );
  HS65_GS_FA1X4 U539 ( .A0(\mul_b1/fa1_c1_r[19] ), .B0(\mul_b1/fa1_c2_r[19] ), 
        .CI(\mul_b1/fa1_s2_r[20] ), .CO(n473), .S0(n466) );
  HS65_GS_FA1X4 U540 ( .A0(n467), .B0(n466), .CI(n465), .CO(n472), .S0(n462)
         );
  HS65_GSS_XOR2X3 U541 ( .A(\mul_b1/fa1_s1_r[21] ), .B(\mul_b1/fa1_s0_r[21] ), 
        .Z(n475) );
  HS65_GS_AND2X4 U542 ( .A(\mul_b1/fa1_s1_r[20] ), .B(\mul_b1/fa1_s0_r[20] ), 
        .Z(n474) );
  HS65_GSS_XNOR2X3 U543 ( .A(n469), .B(n468), .Z(n1777) );
  HS65_GS_NOR2X2 U544 ( .A(n1778), .B(n1777), .Z(n1776) );
  HS65_GS_NOR2X2 U545 ( .A(n470), .B(n1776), .Z(n1126) );
  HS65_GS_FA1X4 U546 ( .A0(n473), .B0(n472), .CI(n471), .CO(n1127), .S0(n1778)
         );
  HS65_GS_FA1X4 U547 ( .A0(\mul_b1/fa1_c1_r[20] ), .B0(\mul_b1/fa1_c2_r[20] ), 
        .CI(\mul_b1/fa1_s2_r[21] ), .CO(n482), .S0(n476) );
  HS65_GS_FA1X4 U548 ( .A0(n476), .B0(n475), .CI(n474), .CO(n481), .S0(n471)
         );
  HS65_GS_FA1X4 U549 ( .A0(n479), .B0(n478), .CI(n477), .CO(n366), .S0(n480)
         );
  HS65_GS_PAO2X4 U550 ( .A(n1126), .B(n1127), .P(n1130), .Z(n1120) );
  HS65_GS_FA1X4 U551 ( .A0(n482), .B0(n481), .CI(n480), .CO(n1121), .S0(n1130)
         );
  HS65_GS_PAO2X4 U552 ( .A(n1125), .B(n1120), .P(n1121), .Z(n1117) );
  HS65_GS_FA1X4 U553 ( .A0(n485), .B0(n484), .CI(n483), .CO(n1114), .S0(n1116)
         );
  HS65_GS_FA1X4 U554 ( .A0(n488), .B0(n487), .CI(n486), .CO(n1110), .S0(n1112)
         );
  HS65_GS_FA1X4 U555 ( .A0(n491), .B0(n490), .CI(n489), .CO(n499), .S0(n497)
         );
  HS65_GS_AND2X4 U556 ( .A(\mul_b1/fa1_c2_r[24] ), .B(\mul_b1/fa1_s2_r[25] ), 
        .Z(n496) );
  HS65_GS_FA1X4 U557 ( .A0(n494), .B0(n493), .CI(n492), .CO(n495), .S0(n486)
         );
  HS65_GS_FA1X4 U558 ( .A0(n497), .B0(n496), .CI(n495), .CO(n1105), .S0(n1108)
         );
  HS65_GS_FA1X4 U559 ( .A0(n500), .B0(n499), .CI(n498), .CO(n1097), .S0(n1104)
         );
  HS65_GS_FA1X4 U560 ( .A0(n503), .B0(n502), .CI(n501), .CO(n1093), .S0(n1095)
         );
  HS65_GS_FA1X4 U561 ( .A0(n506), .B0(n505), .CI(n504), .CO(n514), .S0(n512)
         );
  HS65_GS_AND2X4 U562 ( .A(\mul_b1/fa1_c2_r[27] ), .B(\mul_b1/fa1_s2_r[28] ), 
        .Z(n511) );
  HS65_GS_FA1X4 U563 ( .A0(n509), .B0(n508), .CI(n507), .CO(n510), .S0(n501)
         );
  HS65_GS_FA1X4 U564 ( .A0(n512), .B0(n511), .CI(n510), .CO(n1082), .S0(n1091)
         );
  HS65_GS_FA1X4 U565 ( .A0(n515), .B0(n514), .CI(n513), .CO(n1087), .S0(n1081)
         );
  HS65_GS_AND2X4 U566 ( .A(\mul_b1/fa1_s1_r[30] ), .B(\mul_b1/fa1_s0_r[30] ), 
        .Z(n519) );
  HS65_GSS_XOR2X3 U567 ( .A(\mul_b1/fa1_s1_r[31] ), .B(\mul_b1/fa1_s0_r[31] ), 
        .Z(n518) );
  HS65_GS_FA1X4 U568 ( .A0(n517), .B0(\mul_b1/fa1_s2_r[30] ), .CI(n516), .CO(
        n521), .S0(n513) );
  HS65_GSS_XOR2X3 U569 ( .A(n520), .B(n521), .Z(n1085) );
  HS65_GS_AND2X4 U570 ( .A(\mul_b1/fa1_s1_r[31] ), .B(\mul_b1/fa1_s0_r[31] ), 
        .Z(n525) );
  HS65_GS_NAND2X2 U571 ( .A(\mul_b1/fa1_s1_r[32] ), .B(\mul_b1/fa1_s0_r[32] ), 
        .Z(n529) );
  HS65_GS_OA12X4 U572 ( .A(\mul_b1/fa1_s1_r[32] ), .B(\mul_b1/fa1_s0_r[32] ), 
        .C(n529), .Z(n524) );
  HS65_GS_FA1X4 U573 ( .A0(n519), .B0(\mul_b1/fa1_s2_r[31] ), .CI(n518), .CO(
        n522), .S0(n520) );
  HS65_GSS_XOR2X3 U574 ( .A(n523), .B(n522), .Z(n1089) );
  HS65_GS_AND2X4 U575 ( .A(n521), .B(n520), .Z(n1088) );
  HS65_GS_AND2X4 U576 ( .A(n523), .B(n522), .Z(n528) );
  HS65_GS_FA1X4 U577 ( .A0(\mul_b1/fa1_s2_r[32] ), .B0(n525), .CI(n524), .CO(
        n526), .S0(n523) );
  HS65_GSS_XOR2X3 U578 ( .A(\mul_b1/fa1_s1_r[33] ), .B(n526), .Z(n527) );
  HS65_GSS_XNOR2X3 U579 ( .A(n528), .B(n527), .Z(n530) );
  HS65_GSS_XOR3X2 U580 ( .A(n530), .B(\mul_b1/fa1_s0_r[33] ), .C(n529), .Z(
        n531) );
  HS65_GSS_XOR2X3 U581 ( .A(\mul_b1/fa1_s2_r[33] ), .B(n531), .Z(n532) );
  HS65_GSS_XOR2X3 U582 ( .A(n533), .B(n532), .Z(\mul_b1/result_sat[15] ) );
  HS65_GS_IVX2 U583 ( .A(x_z1[15]), .Z(n1365) );
  HS65_GS_BFX4 U584 ( .A(valid_in), .Z(n1366) );
  HS65_GS_BFX4 U585 ( .A(n1366), .Z(n1792) );
  HS65_GS_IVX2 U586 ( .A(y_z1[15]), .Z(n1635) );
  HS65_GS_IVX2 U587 ( .A(y_z1[14]), .Z(n1637) );
  HS65_GS_IVX2 U588 ( .A(y_z1[13]), .Z(n1639) );
  HS65_GS_IVX2 U589 ( .A(y_z1[12]), .Z(n1641) );
  HS65_GS_IVX2 U590 ( .A(y_z1[11]), .Z(n1643) );
  HS65_GS_IVX2 U591 ( .A(y_z1[10]), .Z(n1645) );
  HS65_GS_IVX2 U592 ( .A(y_z1[9]), .Z(n1647) );
  HS65_GS_IVX2 U593 ( .A(y_z1[8]), .Z(n1649) );
  HS65_GS_IVX2 U594 ( .A(y_z1[7]), .Z(n1651) );
  HS65_GS_IVX2 U595 ( .A(y_z1[6]), .Z(n1653) );
  HS65_GS_IVX2 U596 ( .A(y_z1[5]), .Z(n1655) );
  HS65_GS_IVX2 U597 ( .A(y_z1[4]), .Z(n1657) );
  HS65_GS_IVX2 U598 ( .A(y_z1[3]), .Z(n1659) );
  HS65_GS_IVX2 U599 ( .A(y_z1[2]), .Z(n1661) );
  HS65_GS_IVX2 U600 ( .A(y_z1[1]), .Z(n1713) );
  HS65_GS_IVX2 U601 ( .A(y_z1[0]), .Z(n1712) );
  HS65_GS_NOR2X2 U602 ( .A(y_z1[15]), .B(n1633), .Z(n1788) );
  HS65_GSS_XOR2X3 U603 ( .A(\mul_a1/fa1_s1_r[32] ), .B(\mul_a1/fa1_s0_r[32] ), 
        .Z(n535) );
  HS65_GS_AND2X4 U604 ( .A(\mul_a1/fa1_s0_r[31] ), .B(\mul_a1/fa1_s1_r[31] ), 
        .Z(n534) );
  HS65_GS_FA1X4 U605 ( .A0(n535), .B0(\mul_a1/fa1_s2_r[32] ), .CI(n534), .CO(
        n809), .S0(n536) );
  HS65_GSS_XOR2X3 U606 ( .A(\mul_a1/fa1_s0_r[31] ), .B(\mul_a1/fa1_s1_r[31] ), 
        .Z(n803) );
  HS65_GS_AND2X4 U607 ( .A(\mul_a1/fa1_s0_r[30] ), .B(\mul_a1/fa1_s1_r[30] ), 
        .Z(n802) );
  HS65_GS_AND2X4 U608 ( .A(n536), .B(n537), .Z(n807) );
  HS65_GSS_XNOR2X3 U609 ( .A(n537), .B(n536), .Z(n948) );
  HS65_GSS_XOR2X3 U610 ( .A(\mul_a1/fa1_s0_r[29] ), .B(\mul_a1/fa1_s1_r[29] ), 
        .Z(n544) );
  HS65_GS_NAND2X2 U611 ( .A(\mul_a1/fa1_s1_r[28] ), .B(\mul_a1/fa1_s0_r[28] ), 
        .Z(n538) );
  HS65_GSS_XNOR2X3 U612 ( .A(n538), .B(\mul_a1/fa1_s2_r[29] ), .Z(n545) );
  HS65_GS_NAND2X2 U613 ( .A(n544), .B(n545), .Z(n795) );
  HS65_GS_IVX2 U614 ( .A(n795), .Z(n540) );
  HS65_GS_IVX2 U615 ( .A(\mul_a1/fa1_s2_r[29] ), .Z(n539) );
  HS65_GS_NOR2X2 U616 ( .A(n539), .B(n538), .Z(n794) );
  HS65_GS_AND2X4 U617 ( .A(\mul_a1/fa1_s1_r[29] ), .B(\mul_a1/fa1_s0_r[29] ), 
        .Z(n801) );
  HS65_GSS_XOR2X3 U618 ( .A(\mul_a1/fa1_s0_r[30] ), .B(\mul_a1/fa1_s1_r[30] ), 
        .Z(n800) );
  HS65_GS_IVX2 U619 ( .A(n799), .Z(n798) );
  HS65_GS_OAI21X2 U620 ( .A(n540), .B(n794), .C(n799), .Z(n945) );
  HS65_GSS_XOR2X3 U621 ( .A(\mul_a1/fa1_s1_r[28] ), .B(\mul_a1/fa1_s0_r[28] ), 
        .Z(n783) );
  HS65_GS_NAND2X2 U622 ( .A(\mul_a1/fa1_s1_r[27] ), .B(\mul_a1/fa1_s0_r[27] ), 
        .Z(n541) );
  HS65_GSS_XNOR2X3 U623 ( .A(n541), .B(\mul_a1/fa1_s2_r[28] ), .Z(n784) );
  HS65_GS_NAND2X2 U624 ( .A(n783), .B(n784), .Z(n782) );
  HS65_GS_IVX2 U625 ( .A(n782), .Z(n547) );
  HS65_GS_IVX2 U626 ( .A(\mul_a1/fa1_s2_r[28] ), .Z(n542) );
  HS65_GS_NOR2X2 U627 ( .A(n542), .B(n541), .Z(n546) );
  HS65_GS_IVX2 U628 ( .A(n546), .Z(n543) );
  HS65_GS_NAND2X2 U629 ( .A(n543), .B(n782), .Z(n793) );
  HS65_GS_OAI21X2 U630 ( .A(n545), .B(n544), .C(n795), .Z(n792) );
  HS65_GS_NAND2X2 U631 ( .A(n793), .B(n792), .Z(n791) );
  HS65_GS_OAI21X2 U632 ( .A(n547), .B(n546), .C(n791), .Z(n954) );
  HS65_GS_NAND2X2 U633 ( .A(\mul_a1/fa1_s2_r[26] ), .B(\mul_a1/fa1_c1_r[25] ), 
        .Z(n550) );
  HS65_GS_IVX2 U634 ( .A(n550), .Z(n552) );
  HS65_GSS_XOR2X3 U635 ( .A(\mul_a1/fa1_s1_r[26] ), .B(\mul_a1/fa1_s0_r[26] ), 
        .Z(n769) );
  HS65_GS_AND2X4 U636 ( .A(\mul_a1/fa1_s0_r[25] ), .B(\mul_a1/fa1_s1_r[25] ), 
        .Z(n548) );
  HS65_GSS_XOR3X2 U637 ( .A(\mul_a1/fa1_s2_r[26] ), .B(\mul_a1/fa1_c1_r[25] ), 
        .C(n548), .Z(n770) );
  HS65_GS_NAND2X2 U638 ( .A(n769), .B(n770), .Z(n768) );
  HS65_GS_IVX2 U639 ( .A(n768), .Z(n551) );
  HS65_GS_OAI21X2 U640 ( .A(\mul_a1/fa1_s2_r[26] ), .B(\mul_a1/fa1_c1_r[25] ), 
        .C(n548), .Z(n549) );
  HS65_GS_AND3X4 U641 ( .A(n768), .B(n550), .C(n549), .Z(n555) );
  HS65_GS_AOI12X2 U642 ( .A(n552), .B(n551), .C(n555), .Z(n778) );
  HS65_GS_NAND2X2 U643 ( .A(\mul_a1/fa1_s1_r[26] ), .B(\mul_a1/fa1_s0_r[26] ), 
        .Z(n779) );
  HS65_GS_IVX2 U644 ( .A(\mul_a1/fa1_s2_r[27] ), .Z(n780) );
  HS65_GSS_XOR2X3 U645 ( .A(n779), .B(n780), .Z(n554) );
  HS65_GSS_XOR2X3 U646 ( .A(\mul_a1/fa1_s1_r[27] ), .B(\mul_a1/fa1_s0_r[27] ), 
        .Z(n553) );
  HS65_GS_NAND2X2 U647 ( .A(n553), .B(n554), .Z(n787) );
  HS65_GS_OAI21X2 U648 ( .A(n554), .B(n553), .C(n787), .Z(n777) );
  HS65_GS_AO12X4 U649 ( .A(n778), .B(n777), .C(n555), .Z(n1434) );
  HS65_GS_NAND2X2 U650 ( .A(\mul_a1/fa1_s2_r[24] ), .B(\mul_a1/fa1_c1_r[23] ), 
        .Z(n558) );
  HS65_GS_IVX2 U651 ( .A(n558), .Z(n560) );
  HS65_GSS_XOR2X3 U652 ( .A(\mul_a1/fa1_s1_r[24] ), .B(\mul_a1/fa1_s0_r[24] ), 
        .Z(n570) );
  HS65_GS_AND2X4 U653 ( .A(\mul_a1/fa1_s0_r[23] ), .B(\mul_a1/fa1_s1_r[23] ), 
        .Z(n556) );
  HS65_GSS_XOR3X2 U654 ( .A(\mul_a1/fa1_s2_r[24] ), .B(\mul_a1/fa1_c1_r[23] ), 
        .C(n556), .Z(n571) );
  HS65_GS_NAND2X2 U655 ( .A(n570), .B(n571), .Z(n569) );
  HS65_GS_IVX2 U656 ( .A(n569), .Z(n559) );
  HS65_GS_OAI21X2 U657 ( .A(\mul_a1/fa1_s2_r[24] ), .B(\mul_a1/fa1_c1_r[23] ), 
        .C(n556), .Z(n557) );
  HS65_GS_AND3X4 U658 ( .A(n569), .B(n558), .C(n557), .Z(n563) );
  HS65_GS_AOI12X2 U659 ( .A(n560), .B(n559), .C(n563), .Z(n575) );
  HS65_GS_NAND2X2 U660 ( .A(\mul_a1/fa1_s1_r[24] ), .B(\mul_a1/fa1_s0_r[24] ), 
        .Z(n763) );
  HS65_GS_IVX2 U661 ( .A(\mul_a1/fa1_s2_r[25] ), .Z(n764) );
  HS65_GSS_XOR3X2 U662 ( .A(n763), .B(\mul_a1/fa1_c1_r[24] ), .C(n764), .Z(
        n562) );
  HS65_GSS_XOR2X3 U663 ( .A(\mul_a1/fa1_s1_r[25] ), .B(\mul_a1/fa1_s0_r[25] ), 
        .Z(n561) );
  HS65_GS_NAND2X2 U664 ( .A(n561), .B(n562), .Z(n766) );
  HS65_GS_OAI21X2 U665 ( .A(n562), .B(n561), .C(n766), .Z(n574) );
  HS65_GS_NAND2X2 U666 ( .A(n575), .B(n574), .Z(n573) );
  HS65_GS_NOR2AX3 U667 ( .A(n573), .B(n563), .Z(n761) );
  HS65_GS_NAND2X2 U668 ( .A(\mul_a1/fa1_s2_r[23] ), .B(\mul_a1/fa1_c1_r[22] ), 
        .Z(n566) );
  HS65_GS_IVX2 U669 ( .A(n566), .Z(n568) );
  HS65_GSS_XOR2X3 U670 ( .A(\mul_a1/fa1_s0_r[23] ), .B(\mul_a1/fa1_s1_r[23] ), 
        .Z(n582) );
  HS65_GS_AND2X4 U671 ( .A(\mul_a1/fa1_s1_r[22] ), .B(\mul_a1/fa1_s0_r[22] ), 
        .Z(n564) );
  HS65_GSS_XOR3X2 U672 ( .A(\mul_a1/fa1_s2_r[23] ), .B(\mul_a1/fa1_c1_r[22] ), 
        .C(n564), .Z(n583) );
  HS65_GS_NAND2X2 U673 ( .A(n582), .B(n583), .Z(n581) );
  HS65_GS_IVX2 U674 ( .A(n581), .Z(n567) );
  HS65_GS_OAI21X2 U675 ( .A(\mul_a1/fa1_s2_r[23] ), .B(\mul_a1/fa1_c1_r[22] ), 
        .C(n564), .Z(n565) );
  HS65_GS_AND3X4 U676 ( .A(n581), .B(n566), .C(n565), .Z(n572) );
  HS65_GS_AOI12X2 U677 ( .A(n568), .B(n567), .C(n572), .Z(n760) );
  HS65_GS_OAI21X2 U678 ( .A(n571), .B(n570), .C(n569), .Z(n759) );
  HS65_GS_NAND2X2 U679 ( .A(n760), .B(n759), .Z(n758) );
  HS65_GS_NOR2AX3 U680 ( .A(n758), .B(n572), .Z(n1438) );
  HS65_GS_OAI21X2 U681 ( .A(n575), .B(n574), .C(n573), .Z(n1437) );
  HS65_GS_NAND2X2 U682 ( .A(\mul_a1/fa1_s2_r[22] ), .B(\mul_a1/fa1_c1_r[21] ), 
        .Z(n578) );
  HS65_GS_IVX2 U683 ( .A(n578), .Z(n580) );
  HS65_GSS_XOR2X3 U684 ( .A(\mul_a1/fa1_s1_r[22] ), .B(\mul_a1/fa1_s0_r[22] ), 
        .Z(n745) );
  HS65_GS_AND2X4 U685 ( .A(\mul_a1/fa1_s1_r[21] ), .B(\mul_a1/fa1_s0_r[21] ), 
        .Z(n576) );
  HS65_GSS_XOR3X2 U686 ( .A(\mul_a1/fa1_s2_r[22] ), .B(\mul_a1/fa1_c1_r[21] ), 
        .C(n576), .Z(n746) );
  HS65_GS_NAND2X2 U687 ( .A(n745), .B(n746), .Z(n744) );
  HS65_GS_IVX2 U688 ( .A(n744), .Z(n579) );
  HS65_GS_OAI21X2 U689 ( .A(\mul_a1/fa1_s2_r[22] ), .B(\mul_a1/fa1_c1_r[21] ), 
        .C(n576), .Z(n577) );
  HS65_GS_AND3X4 U690 ( .A(n744), .B(n578), .C(n577), .Z(n584) );
  HS65_GS_AOI12X2 U691 ( .A(n580), .B(n579), .C(n584), .Z(n757) );
  HS65_GS_OAI21X2 U692 ( .A(n583), .B(n582), .C(n581), .Z(n756) );
  HS65_GS_NAND2X2 U693 ( .A(n757), .B(n756), .Z(n755) );
  HS65_GS_NOR2AX3 U694 ( .A(n755), .B(n584), .Z(n1442) );
  HS65_GS_AND2X4 U695 ( .A(\mul_a1/fa1_s2_r[14] ), .B(\mul_a1/fa1_c1_r[13] ), 
        .Z(n587) );
  HS65_GSS_XOR3X2 U696 ( .A(\mul_a1/fa1_s1_r[15] ), .B(\mul_a1/fa1_c0_r[14] ), 
        .C(\mul_a1/fa1_s0_r[15] ), .Z(n649) );
  HS65_GSS_XOR3X2 U697 ( .A(n649), .B(\mul_a1/fa1_c1_r[14] ), .C(
        \mul_a1/fa1_s2_r[15] ), .Z(n651) );
  HS65_GSS_XOR2X3 U698 ( .A(n651), .B(n650), .Z(n586) );
  HS65_GSS_XOR2X3 U699 ( .A(\mul_a1/fa1_s2_r[14] ), .B(\mul_a1/fa1_c1_r[13] ), 
        .Z(n639) );
  HS65_GS_FA1X4 U700 ( .A0(\mul_a1/fa1_s0_r[14] ), .B0(\mul_a1/fa1_s1_r[14] ), 
        .CI(\mul_a1/fa1_c0_r[13] ), .CO(n650), .S0(n638) );
  HS65_GS_FA1X4 U701 ( .A0(n587), .B0(n586), .CI(n585), .CO(n657), .S0(n647)
         );
  HS65_GS_AND2X4 U702 ( .A(\mul_a1/fa1_c1_r[11] ), .B(\mul_a1/fa1_s2_r[12] ), 
        .Z(n589) );
  HS65_GSS_XOR2X3 U703 ( .A(\mul_a1/fa1_c1_r[11] ), .B(\mul_a1/fa1_s2_r[12] ), 
        .Z(n594) );
  HS65_GS_PAO2X4 U704 ( .A(\mul_a1/fa1_s1_r[11] ), .B(\mul_a1/fa1_s0_r[11] ), 
        .P(\mul_a1/fa1_c0_r[10] ), .Z(n593) );
  HS65_GS_PAO2X4 U705 ( .A(n595), .B(n594), .P(n593), .Z(n590) );
  HS65_GS_NOR2X2 U706 ( .A(n589), .B(n590), .Z(n592) );
  HS65_GS_FA1X4 U707 ( .A0(\mul_a1/fa1_s0_r[12] ), .B0(\mul_a1/fa1_s1_r[12] ), 
        .CI(\mul_a1/fa1_c0_r[11] ), .CO(n642), .S0(n595) );
  HS65_GS_FA1X4 U708 ( .A0(\mul_a1/fa1_s0_r[13] ), .B0(\mul_a1/fa1_s1_r[13] ), 
        .CI(\mul_a1/fa1_c0_r[12] ), .CO(n637), .S0(n641) );
  HS65_GSS_XOR2X3 U709 ( .A(\mul_a1/fa1_s2_r[13] ), .B(\mul_a1/fa1_c1_r[12] ), 
        .Z(n640) );
  HS65_GS_NAND3X2 U710 ( .A(n593), .B(n595), .C(n589), .Z(n588) );
  HS65_GS_OAI21X2 U711 ( .A(n590), .B(n589), .C(n588), .Z(n630) );
  HS65_GS_NOR2X2 U712 ( .A(n632), .B(n630), .Z(n591) );
  HS65_GS_NOR2X2 U713 ( .A(n592), .B(n591), .Z(n636) );
  HS65_GSS_XOR3X2 U714 ( .A(n595), .B(n594), .C(n593), .Z(n629) );
  HS65_GSS_XNOR3X2 U715 ( .A(\mul_a1/fa1_s1_r[11] ), .B(\mul_a1/fa1_s0_r[11] ), 
        .C(\mul_a1/fa1_c0_r[10] ), .Z(n620) );
  HS65_GS_PAOI2X1 U716 ( .A(\mul_a1/fa1_s1_r[10] ), .B(\mul_a1/fa1_c0_r[9] ), 
        .P(\mul_a1/fa1_s0_r[10] ), .Z(n621) );
  HS65_GS_NOR2X2 U717 ( .A(n620), .B(n621), .Z(n628) );
  HS65_GSS_XNOR3X2 U718 ( .A(\mul_a1/fa1_c0_r[8] ), .B(\mul_a1/fa1_s1_r[9] ), 
        .C(\mul_a1/fa1_s0_r[9] ), .Z(n613) );
  HS65_GS_NAND2X2 U719 ( .A(\mul_a1/fa1_c0_r[7] ), .B(\mul_a1/fa1_s0_r[8] ), 
        .Z(n596) );
  HS65_GS_NOR2X2 U720 ( .A(n613), .B(n596), .Z(n619) );
  HS65_GS_PAOI2X1 U721 ( .A(\mul_a1/fa1_c0_r[8] ), .B(\mul_a1/fa1_s1_r[9] ), 
        .P(\mul_a1/fa1_s0_r[9] ), .Z(n622) );
  HS65_GSS_XNOR3X2 U722 ( .A(\mul_a1/fa1_s1_r[10] ), .B(\mul_a1/fa1_c0_r[9] ), 
        .C(\mul_a1/fa1_s0_r[10] ), .Z(n623) );
  HS65_GSS_XOR2X3 U723 ( .A(n622), .B(n623), .Z(n618) );
  HS65_GSS_XNOR2X3 U724 ( .A(\mul_a1/fa1_c0_r[6] ), .B(\mul_a1/fa1_s0_r[7] ), 
        .Z(n604) );
  HS65_GS_NAND2X2 U725 ( .A(\mul_a1/fa1_c0_r[5] ), .B(\mul_a1/fa1_s0_r[6] ), 
        .Z(n597) );
  HS65_GS_NOR2X2 U726 ( .A(n604), .B(n597), .Z(n610) );
  HS65_GSS_XNOR2X3 U727 ( .A(\mul_a1/fa1_c0_r[7] ), .B(\mul_a1/fa1_s0_r[8] ), 
        .Z(n612) );
  HS65_GS_IVX2 U728 ( .A(n612), .Z(n609) );
  HS65_GSS_XNOR2X3 U729 ( .A(\mul_a1/fa1_c0_r[4] ), .B(\mul_a1/fa1_s0_r[5] ), 
        .Z(n599) );
  HS65_GS_NAND2X2 U730 ( .A(\mul_a1/fa1_c0_r[3] ), .B(\mul_a1/fa1_s0_r[4] ), 
        .Z(n598) );
  HS65_GS_NOR2X2 U731 ( .A(n599), .B(n598), .Z(n601) );
  HS65_GSS_XNOR2X3 U732 ( .A(\mul_a1/fa1_c0_r[5] ), .B(\mul_a1/fa1_s0_r[6] ), 
        .Z(n603) );
  HS65_GS_IVX2 U733 ( .A(n603), .Z(n600) );
  HS65_GS_AND2X4 U734 ( .A(n601), .B(n600), .Z(n607) );
  HS65_GS_NAND2X2 U735 ( .A(\mul_a1/fa1_c0_r[4] ), .B(\mul_a1/fa1_s0_r[5] ), 
        .Z(n602) );
  HS65_GS_NOR2X2 U736 ( .A(n603), .B(n602), .Z(n606) );
  HS65_GS_IVX2 U737 ( .A(n604), .Z(n605) );
  HS65_GS_PAO2X4 U738 ( .A(n607), .B(n606), .P(n605), .Z(n608) );
  HS65_GS_PAO2X4 U739 ( .A(n610), .B(n609), .P(n608), .Z(n616) );
  HS65_GS_NAND2X2 U740 ( .A(\mul_a1/fa1_c0_r[6] ), .B(\mul_a1/fa1_s0_r[7] ), 
        .Z(n611) );
  HS65_GS_NOR2X2 U741 ( .A(n612), .B(n611), .Z(n615) );
  HS65_GS_IVX2 U742 ( .A(n613), .Z(n614) );
  HS65_GS_PAO2X4 U743 ( .A(n616), .B(n615), .P(n614), .Z(n617) );
  HS65_GS_PAO2X4 U744 ( .A(n619), .B(n618), .P(n617), .Z(n626) );
  HS65_GSS_XOR2X3 U745 ( .A(n621), .B(n620), .Z(n625) );
  HS65_GS_NOR2X2 U746 ( .A(n623), .B(n622), .Z(n624) );
  HS65_GS_PAO2X4 U747 ( .A(n626), .B(n625), .P(n624), .Z(n627) );
  HS65_GS_PAOI2X1 U748 ( .A(n629), .B(n628), .P(n627), .Z(n634) );
  HS65_GS_IVX2 U749 ( .A(n630), .Z(n631) );
  HS65_GS_NOR2X2 U750 ( .A(n632), .B(n631), .Z(n633) );
  HS65_GS_NOR2X2 U751 ( .A(n634), .B(n633), .Z(n635) );
  HS65_GS_NOR2X2 U752 ( .A(n636), .B(n635), .Z(n1730) );
  HS65_GS_AND2X4 U753 ( .A(\mul_a1/fa1_s2_r[13] ), .B(\mul_a1/fa1_c1_r[12] ), 
        .Z(n645) );
  HS65_GS_FA1X4 U754 ( .A0(n639), .B0(n638), .CI(n637), .CO(n585), .S0(n644)
         );
  HS65_GS_FA1X4 U755 ( .A0(n642), .B0(n641), .CI(n640), .CO(n643), .S0(n632)
         );
  HS65_GS_NOR2X2 U756 ( .A(n1731), .B(n1730), .Z(n1729) );
  HS65_GS_NOR2X2 U757 ( .A(n1730), .B(n1729), .Z(n646) );
  HS65_GS_NAND2X2 U758 ( .A(n647), .B(n646), .Z(n648) );
  HS65_GS_FA1X4 U759 ( .A0(n645), .B0(n644), .CI(n643), .CO(n1452), .S0(n1731)
         );
  HS65_GSS_XOR2X3 U760 ( .A(n647), .B(n646), .Z(n1451) );
  HS65_GS_NAND2X2 U761 ( .A(n1452), .B(n1451), .Z(n1450) );
  HS65_GS_NAND2X2 U762 ( .A(n648), .B(n1450), .Z(n656) );
  HS65_GS_AND2X4 U763 ( .A(n657), .B(n656), .Z(n659) );
  HS65_GS_AND2X4 U764 ( .A(\mul_a1/fa1_c1_r[14] ), .B(\mul_a1/fa1_s2_r[15] ), 
        .Z(n652) );
  HS65_GS_CB4I6X4 U765 ( .A(\mul_a1/fa1_c1_r[14] ), .B(\mul_a1/fa1_s2_r[15] ), 
        .C(n649), .D(n652), .Z(n663) );
  HS65_GS_IVX2 U766 ( .A(n663), .Z(n653) );
  HS65_GS_AND2X4 U767 ( .A(n651), .B(n650), .Z(n664) );
  HS65_GS_MUXI21X2 U768 ( .D0(n653), .D1(n652), .S0(n664), .Z(n661) );
  HS65_GS_PAOI2X1 U769 ( .A(\mul_a1/fa1_s1_r[15] ), .B(\mul_a1/fa1_c0_r[14] ), 
        .P(\mul_a1/fa1_s0_r[15] ), .Z(n667) );
  HS65_GS_IVX2 U770 ( .A(\mul_a1/fa1_s2_r[16] ), .Z(n668) );
  HS65_GSS_XOR3X2 U771 ( .A(n667), .B(\mul_a1/fa1_c1_r[15] ), .C(n668), .Z(
        n655) );
  HS65_GSS_XOR3X2 U772 ( .A(\mul_a1/fa1_s1_r[16] ), .B(\mul_a1/fa1_c0_r[15] ), 
        .C(\mul_a1/fa1_s0_r[16] ), .Z(n654) );
  HS65_GS_NAND2X2 U773 ( .A(n654), .B(n655), .Z(n670) );
  HS65_GS_OAI21X2 U774 ( .A(n655), .B(n654), .C(n670), .Z(n660) );
  HS65_GSS_XOR2X3 U775 ( .A(n661), .B(n660), .Z(n979) );
  HS65_GSS_XNOR2X3 U776 ( .A(n657), .B(n656), .Z(n980) );
  HS65_GS_NOR2X2 U777 ( .A(n979), .B(n980), .Z(n658) );
  HS65_GS_NOR2X2 U778 ( .A(n659), .B(n658), .Z(n665) );
  HS65_GS_NAND2X2 U779 ( .A(n661), .B(n660), .Z(n662) );
  HS65_GS_OAI21X2 U780 ( .A(n664), .B(n663), .C(n662), .Z(n666) );
  HS65_GS_NAND2X2 U781 ( .A(n665), .B(n666), .Z(n674) );
  HS65_GSS_XOR2X3 U782 ( .A(n666), .B(n665), .Z(n1735) );
  HS65_GS_IVX2 U783 ( .A(\mul_a1/fa1_c1_r[15] ), .Z(n669) );
  HS65_GS_NAND2X2 U784 ( .A(\mul_a1/fa1_c1_r[15] ), .B(\mul_a1/fa1_s2_r[16] ), 
        .Z(n671) );
  HS65_GS_CBI4I1X3 U785 ( .A(n669), .B(n668), .C(n667), .D(n671), .Z(n678) );
  HS65_GS_IVX2 U786 ( .A(n670), .Z(n679) );
  HS65_GS_MUX21X4 U787 ( .D0(n678), .D1(n671), .S0(n679), .Z(n676) );
  HS65_GS_PAOI2X1 U788 ( .A(\mul_a1/fa1_s1_r[16] ), .B(\mul_a1/fa1_c0_r[15] ), 
        .P(\mul_a1/fa1_s0_r[16] ), .Z(n680) );
  HS65_GS_IVX2 U789 ( .A(\mul_a1/fa1_s2_r[17] ), .Z(n681) );
  HS65_GSS_XOR3X2 U790 ( .A(n680), .B(\mul_a1/fa1_c1_r[16] ), .C(n681), .Z(
        n673) );
  HS65_GSS_XOR3X2 U791 ( .A(\mul_a1/fa1_s1_r[17] ), .B(\mul_a1/fa1_c0_r[16] ), 
        .C(\mul_a1/fa1_s0_r[17] ), .Z(n672) );
  HS65_GS_NAND2X2 U792 ( .A(n672), .B(n673), .Z(n683) );
  HS65_GS_OAI21X2 U793 ( .A(n673), .B(n672), .C(n683), .Z(n675) );
  HS65_GSS_XOR2X3 U794 ( .A(n676), .B(n675), .Z(n1734) );
  HS65_GS_NAND2X2 U795 ( .A(n1735), .B(n1734), .Z(n1733) );
  HS65_GS_NAND2X2 U796 ( .A(n674), .B(n1733), .Z(n688) );
  HS65_GS_NAND2X2 U797 ( .A(n676), .B(n675), .Z(n677) );
  HS65_GS_OAI21X2 U798 ( .A(n679), .B(n678), .C(n677), .Z(n687) );
  HS65_GS_NOR2X2 U799 ( .A(n688), .B(n687), .Z(n690) );
  HS65_GS_IVX2 U800 ( .A(\mul_a1/fa1_c1_r[16] ), .Z(n682) );
  HS65_GS_NAND2X2 U801 ( .A(\mul_a1/fa1_c1_r[16] ), .B(\mul_a1/fa1_s2_r[17] ), 
        .Z(n684) );
  HS65_GS_CBI4I1X3 U802 ( .A(n682), .B(n681), .C(n680), .D(n684), .Z(n694) );
  HS65_GS_IVX2 U803 ( .A(n683), .Z(n695) );
  HS65_GS_MUX21X4 U804 ( .D0(n694), .D1(n684), .S0(n695), .Z(n692) );
  HS65_GS_PAOI2X1 U805 ( .A(\mul_a1/fa1_s1_r[17] ), .B(\mul_a1/fa1_c0_r[16] ), 
        .P(\mul_a1/fa1_s0_r[17] ), .Z(n696) );
  HS65_GS_IVX2 U806 ( .A(\mul_a1/fa1_s2_r[18] ), .Z(n697) );
  HS65_GSS_XOR3X2 U807 ( .A(n696), .B(\mul_a1/fa1_c1_r[17] ), .C(n697), .Z(
        n686) );
  HS65_GSS_XOR3X2 U808 ( .A(\mul_a1/fa1_s1_r[18] ), .B(\mul_a1/fa1_c0_r[17] ), 
        .C(\mul_a1/fa1_s0_r[18] ), .Z(n685) );
  HS65_GS_NAND2X2 U809 ( .A(n685), .B(n686), .Z(n699) );
  HS65_GS_OAI21X2 U810 ( .A(n686), .B(n685), .C(n699), .Z(n691) );
  HS65_GSS_XOR2X3 U811 ( .A(n692), .B(n691), .Z(n976) );
  HS65_GSS_XNOR2X3 U812 ( .A(n688), .B(n687), .Z(n977) );
  HS65_GS_NOR2X2 U813 ( .A(n976), .B(n977), .Z(n689) );
  HS65_GS_NOR2X2 U814 ( .A(n690), .B(n689), .Z(n704) );
  HS65_GS_NAND2X2 U815 ( .A(n692), .B(n691), .Z(n693) );
  HS65_GS_OAI21X2 U816 ( .A(n695), .B(n694), .C(n693), .Z(n703) );
  HS65_GS_NOR2X2 U817 ( .A(n704), .B(n703), .Z(n706) );
  HS65_GS_IVX2 U818 ( .A(\mul_a1/fa1_c1_r[17] ), .Z(n698) );
  HS65_GS_NAND2X2 U819 ( .A(\mul_a1/fa1_c1_r[17] ), .B(\mul_a1/fa1_s2_r[18] ), 
        .Z(n700) );
  HS65_GS_CBI4I1X3 U820 ( .A(n698), .B(n697), .C(n696), .D(n700), .Z(n710) );
  HS65_GS_IVX2 U821 ( .A(n699), .Z(n711) );
  HS65_GS_MUX21X4 U822 ( .D0(n710), .D1(n700), .S0(n711), .Z(n708) );
  HS65_GS_PAOI2X1 U823 ( .A(\mul_a1/fa1_s1_r[18] ), .B(\mul_a1/fa1_c0_r[17] ), 
        .P(\mul_a1/fa1_s0_r[18] ), .Z(n714) );
  HS65_GS_IVX2 U824 ( .A(\mul_a1/fa1_s2_r[19] ), .Z(n715) );
  HS65_GSS_XOR3X2 U825 ( .A(n714), .B(\mul_a1/fa1_c1_r[18] ), .C(n715), .Z(
        n702) );
  HS65_GSS_XOR2X3 U826 ( .A(\mul_a1/fa1_s1_r[19] ), .B(\mul_a1/fa1_s0_r[19] ), 
        .Z(n701) );
  HS65_GS_NAND2X2 U827 ( .A(n701), .B(n702), .Z(n717) );
  HS65_GS_OAI21X2 U828 ( .A(n702), .B(n701), .C(n717), .Z(n707) );
  HS65_GSS_XOR2X3 U829 ( .A(n708), .B(n707), .Z(n973) );
  HS65_GSS_XNOR2X3 U830 ( .A(n704), .B(n703), .Z(n974) );
  HS65_GS_NOR2X2 U831 ( .A(n973), .B(n974), .Z(n705) );
  HS65_GS_NOR2X2 U832 ( .A(n706), .B(n705), .Z(n713) );
  HS65_GS_NAND2X2 U833 ( .A(n708), .B(n707), .Z(n709) );
  HS65_GS_OAI21X2 U834 ( .A(n711), .B(n710), .C(n709), .Z(n712) );
  HS65_GS_NAND2X2 U835 ( .A(n713), .B(n712), .Z(n721) );
  HS65_GSS_XOR2X3 U836 ( .A(n713), .B(n712), .Z(n1739) );
  HS65_GS_IVX2 U837 ( .A(\mul_a1/fa1_c1_r[18] ), .Z(n716) );
  HS65_GS_NAND2X2 U838 ( .A(\mul_a1/fa1_c1_r[18] ), .B(\mul_a1/fa1_s2_r[19] ), 
        .Z(n718) );
  HS65_GS_CBI4I1X3 U839 ( .A(n716), .B(n715), .C(n714), .D(n718), .Z(n725) );
  HS65_GS_IVX2 U840 ( .A(n717), .Z(n726) );
  HS65_GS_MUX21X4 U841 ( .D0(n725), .D1(n718), .S0(n726), .Z(n723) );
  HS65_GS_NAND2X2 U842 ( .A(\mul_a1/fa1_s1_r[19] ), .B(\mul_a1/fa1_s0_r[19] ), 
        .Z(n727) );
  HS65_GS_IVX2 U843 ( .A(\mul_a1/fa1_s2_r[20] ), .Z(n728) );
  HS65_GSS_XOR3X2 U844 ( .A(n727), .B(\mul_a1/fa1_c1_r[19] ), .C(n728), .Z(
        n720) );
  HS65_GSS_XOR2X3 U845 ( .A(\mul_a1/fa1_s1_r[20] ), .B(\mul_a1/fa1_s0_r[20] ), 
        .Z(n719) );
  HS65_GS_NAND2X2 U846 ( .A(n719), .B(n720), .Z(n730) );
  HS65_GS_OAI21X2 U847 ( .A(n720), .B(n719), .C(n730), .Z(n722) );
  HS65_GSS_XOR2X3 U848 ( .A(n723), .B(n722), .Z(n1738) );
  HS65_GS_NAND2X2 U849 ( .A(n1739), .B(n1738), .Z(n1737) );
  HS65_GS_NAND2X2 U850 ( .A(n721), .B(n1737), .Z(n735) );
  HS65_GS_NAND2X2 U851 ( .A(n723), .B(n722), .Z(n724) );
  HS65_GS_OAI21X2 U852 ( .A(n726), .B(n725), .C(n724), .Z(n734) );
  HS65_GS_NOR2X2 U853 ( .A(n735), .B(n734), .Z(n737) );
  HS65_GS_IVX2 U854 ( .A(\mul_a1/fa1_c1_r[19] ), .Z(n729) );
  HS65_GS_NAND2X2 U855 ( .A(\mul_a1/fa1_c1_r[19] ), .B(\mul_a1/fa1_s2_r[20] ), 
        .Z(n731) );
  HS65_GS_CBI4I1X3 U856 ( .A(n729), .B(n728), .C(n727), .D(n731), .Z(n750) );
  HS65_GS_IVX2 U857 ( .A(n730), .Z(n751) );
  HS65_GS_MUX21X4 U858 ( .D0(n750), .D1(n731), .S0(n751), .Z(n748) );
  HS65_GS_AND2X4 U859 ( .A(\mul_a1/fa1_s0_r[20] ), .B(\mul_a1/fa1_s1_r[20] ), 
        .Z(n738) );
  HS65_GSS_XOR3X2 U860 ( .A(\mul_a1/fa1_s2_r[21] ), .B(\mul_a1/fa1_c1_r[20] ), 
        .C(n738), .Z(n733) );
  HS65_GSS_XOR2X3 U861 ( .A(\mul_a1/fa1_s1_r[21] ), .B(\mul_a1/fa1_s0_r[21] ), 
        .Z(n732) );
  HS65_GS_NAND2X2 U862 ( .A(n732), .B(n733), .Z(n741) );
  HS65_GS_OAI21X2 U863 ( .A(n733), .B(n732), .C(n741), .Z(n747) );
  HS65_GSS_XOR2X3 U864 ( .A(n748), .B(n747), .Z(n970) );
  HS65_GSS_XNOR2X3 U865 ( .A(n735), .B(n734), .Z(n971) );
  HS65_GS_NOR2X2 U866 ( .A(n970), .B(n971), .Z(n736) );
  HS65_GS_NOR2X2 U867 ( .A(n737), .B(n736), .Z(n965) );
  HS65_GS_NAND2X2 U868 ( .A(\mul_a1/fa1_s2_r[21] ), .B(\mul_a1/fa1_c1_r[20] ), 
        .Z(n740) );
  HS65_GS_IVX2 U869 ( .A(n740), .Z(n743) );
  HS65_GS_IVX2 U870 ( .A(n741), .Z(n742) );
  HS65_GS_OAI21X2 U871 ( .A(\mul_a1/fa1_s2_r[21] ), .B(\mul_a1/fa1_c1_r[20] ), 
        .C(n738), .Z(n739) );
  HS65_GS_AND3X4 U872 ( .A(n741), .B(n740), .C(n739), .Z(n752) );
  HS65_GS_AOI12X2 U873 ( .A(n743), .B(n742), .C(n752), .Z(n754) );
  HS65_GS_OAI21X2 U874 ( .A(n746), .B(n745), .C(n744), .Z(n753) );
  HS65_GSS_XOR2X3 U875 ( .A(n754), .B(n753), .Z(n967) );
  HS65_GS_NAND2X2 U876 ( .A(n748), .B(n747), .Z(n749) );
  HS65_GS_OAI21X2 U877 ( .A(n751), .B(n750), .C(n749), .Z(n964) );
  HS65_GS_PAOI2X1 U878 ( .A(n965), .B(n967), .P(n964), .Z(n1446) );
  HS65_GS_AOI12X2 U879 ( .A(n754), .B(n753), .C(n752), .Z(n1445) );
  HS65_GS_OAI21X2 U880 ( .A(n757), .B(n756), .C(n755), .Z(n1444) );
  HS65_GS_OAI21X2 U881 ( .A(n760), .B(n759), .C(n758), .Z(n1440) );
  HS65_GS_NOR2X2 U882 ( .A(n761), .B(n762), .Z(n771) );
  HS65_GSS_XNOR2X3 U883 ( .A(n762), .B(n761), .Z(n1743) );
  HS65_GS_IVX2 U884 ( .A(\mul_a1/fa1_c1_r[24] ), .Z(n765) );
  HS65_GS_NAND2X2 U885 ( .A(\mul_a1/fa1_c1_r[24] ), .B(\mul_a1/fa1_s2_r[25] ), 
        .Z(n767) );
  HS65_GS_CBI4I1X3 U886 ( .A(n765), .B(n764), .C(n763), .D(n767), .Z(n775) );
  HS65_GS_IVX2 U887 ( .A(n766), .Z(n776) );
  HS65_GS_MUX21X4 U888 ( .D0(n775), .D1(n767), .S0(n776), .Z(n773) );
  HS65_GS_OAI21X2 U889 ( .A(n770), .B(n769), .C(n768), .Z(n772) );
  HS65_GSS_XNOR2X3 U890 ( .A(n773), .B(n772), .Z(n1742) );
  HS65_GS_NOR2X2 U891 ( .A(n1743), .B(n1742), .Z(n1741) );
  HS65_GS_NOR2X2 U892 ( .A(n771), .B(n1741), .Z(n941) );
  HS65_GS_NAND2X2 U893 ( .A(n773), .B(n772), .Z(n774) );
  HS65_GS_OA12X4 U894 ( .A(n776), .B(n775), .C(n774), .Z(n940) );
  HS65_GSS_XNOR2X3 U895 ( .A(n778), .B(n777), .Z(n942) );
  HS65_GS_PAOI2X1 U896 ( .A(n941), .B(n940), .P(n942), .Z(n1433) );
  HS65_GS_NOR2X2 U897 ( .A(n780), .B(n779), .Z(n789) );
  HS65_GS_IVX2 U898 ( .A(n789), .Z(n781) );
  HS65_GS_NAND2X2 U899 ( .A(n781), .B(n787), .Z(n786) );
  HS65_GS_OAI21X2 U900 ( .A(n784), .B(n783), .C(n782), .Z(n785) );
  HS65_GS_NAND2X2 U901 ( .A(n786), .B(n785), .Z(n788) );
  HS65_GS_OA12X4 U902 ( .A(n786), .B(n785), .C(n788), .Z(n1432) );
  HS65_GS_IVX2 U903 ( .A(n787), .Z(n790) );
  HS65_GS_OAI21X2 U904 ( .A(n790), .B(n789), .C(n788), .Z(n950) );
  HS65_GS_OA12X4 U905 ( .A(n793), .B(n792), .C(n791), .Z(n949) );
  HS65_GS_IVX2 U906 ( .A(n794), .Z(n796) );
  HS65_GS_NAND2X2 U907 ( .A(n796), .B(n795), .Z(n797) );
  HS65_GS_MUXI21X2 U908 ( .D0(n799), .D1(n798), .S0(n797), .Z(n952) );
  HS65_GS_FA1X4 U909 ( .A0(n801), .B0(n800), .CI(\mul_a1/fa1_s2_r[30] ), .CO(
        n804), .S0(n799) );
  HS65_GS_FA1X4 U910 ( .A0(\mul_a1/fa1_s2_r[31] ), .B0(n803), .CI(n802), .CO(
        n537), .S0(n805) );
  HS65_GSS_XNOR2X3 U911 ( .A(n804), .B(n805), .Z(n943) );
  HS65_GS_NAND2X2 U912 ( .A(n805), .B(n804), .Z(n946) );
  HS65_GSS_XOR2X3 U913 ( .A(n807), .B(n806), .Z(n808) );
  HS65_GSS_XNOR2X3 U914 ( .A(n809), .B(n808), .Z(n812) );
  HS65_GS_NAND2X2 U915 ( .A(\mul_a1/fa1_s1_r[32] ), .B(\mul_a1/fa1_s0_r[32] ), 
        .Z(n810) );
  HS65_GSS_XNOR3X2 U916 ( .A(n810), .B(\mul_a1/fa1_s0_r[33] ), .C(
        \mul_a1/fa1_s1_r[33] ), .Z(n811) );
  HS65_GSS_XOR3X2 U917 ( .A(\mul_a1/fa1_s2_r[33] ), .B(n812), .C(n811), .Z(
        \mul_a1/result_sat[15] ) );
  HS65_GS_IVX2 U918 ( .A(y_z2[15]), .Z(n1710) );
  HS65_GS_HA1X4 U919 ( .A0(n1713), .B0(n1712), .CO(n1400) );
  HS65_GS_NOR2X2 U920 ( .A(y_z1[15]), .B(n1431), .Z(n1632) );
  HS65_GSS_XNOR2X6 U921 ( .A(n1632), .B(n1635), .Z(\mul_a1/fa1_s0[29] ) );
  HS65_GS_IVX2 U922 ( .A(x_reg2[0]), .Z(n1677) );
  HS65_GS_IVX2 U923 ( .A(x_reg2[2]), .Z(n1715) );
  HS65_GS_NOR2X2 U924 ( .A(n1677), .B(n1715), .Z(\mul_b2/fa1_c0[4] ) );
  HS65_GS_IVX2 U925 ( .A(x_reg2[15]), .Z(n1727) );
  HS65_GS_IVX2 U926 ( .A(x_reg2[14]), .Z(n1728) );
  HS65_GS_IVX2 U927 ( .A(x_reg2[13]), .Z(n1726) );
  HS65_GS_IVX2 U928 ( .A(x_reg2[12]), .Z(n1725) );
  HS65_GS_IVX2 U929 ( .A(x_reg2[11]), .Z(n1724) );
  HS65_GS_IVX2 U930 ( .A(x_reg2[10]), .Z(n1723) );
  HS65_GS_IVX2 U931 ( .A(x_reg2[9]), .Z(n1722) );
  HS65_GS_IVX2 U932 ( .A(x_reg2[8]), .Z(n1721) );
  HS65_GS_IVX2 U933 ( .A(x_reg2[7]), .Z(n1720) );
  HS65_GS_IVX2 U934 ( .A(x_reg2[6]), .Z(n1719) );
  HS65_GS_IVX2 U935 ( .A(x_reg2[5]), .Z(n1718) );
  HS65_GS_IVX2 U936 ( .A(x_reg2[4]), .Z(n1717) );
  HS65_GS_IVX2 U937 ( .A(x_reg2[3]), .Z(n1716) );
  HS65_GS_IVX2 U938 ( .A(x_reg2[1]), .Z(n1714) );
  HS65_GS_NOR2X3 U939 ( .A(x_reg2[15]), .B(n1662), .Z(n1786) );
  HS65_GS_FA1X4 U940 ( .A0(n815), .B0(n814), .CI(n813), .CO(n822), .S0(n829)
         );
  HS65_GS_FA1X4 U941 ( .A0(n818), .B0(n817), .CI(n816), .CO(n813), .S0(n828)
         );
  HS65_GS_FA1X4 U942 ( .A0(n821), .B0(n820), .CI(n819), .CO(n816), .S0(n827)
         );
  HS65_GS_NOR3X1 U943 ( .A(n829), .B(n828), .C(n827), .Z(n826) );
  HS65_GS_FA1X4 U944 ( .A0(n824), .B0(n823), .CI(n822), .CO(n237), .S0(n825)
         );
  HS65_GS_IVX2 U945 ( .A(n825), .Z(n831) );
  HS65_GS_AOI12X2 U946 ( .A(n826), .B(n831), .C(\mul_b2/result_sat[15] ), .Z(
        n1033) );
  HS65_GS_IVX2 U947 ( .A(n1033), .Z(n868) );
  HS65_GS_NAND3X2 U948 ( .A(n829), .B(n828), .C(n827), .Z(n830) );
  HS65_GS_OAI21X2 U949 ( .A(n831), .B(n830), .C(\mul_b2/result_sat[15] ), .Z(
        n1034) );
  HS65_GS_IVX2 U950 ( .A(n1034), .Z(n1018) );
  HS65_GS_AO112X4 U951 ( .A(n834), .B(n833), .C(n1018), .D(n832), .Z(n835) );
  HS65_GS_NAND2X2 U952 ( .A(n868), .B(n835), .Z(\mul_b2/result_sat[11] ) );
  HS65_GS_AO112X4 U953 ( .A(n838), .B(n837), .C(n1018), .D(n836), .Z(n839) );
  HS65_GS_NAND2X2 U954 ( .A(n868), .B(n839), .Z(\mul_b2/result_sat[10] ) );
  HS65_GS_AO112X4 U955 ( .A(n842), .B(n841), .C(n1018), .D(n840), .Z(n843) );
  HS65_GS_NAND2X2 U956 ( .A(n868), .B(n843), .Z(\mul_b2/result_sat[9] ) );
  HS65_GS_AO112X4 U957 ( .A(n846), .B(n845), .C(n1018), .D(n844), .Z(n847) );
  HS65_GS_NAND2X2 U958 ( .A(n868), .B(n847), .Z(\mul_b2/result_sat[8] ) );
  HS65_GS_AO112X4 U959 ( .A(n850), .B(n849), .C(n1018), .D(n848), .Z(n851) );
  HS65_GS_NAND2X2 U960 ( .A(n868), .B(n851), .Z(\mul_b2/result_sat[7] ) );
  HS65_GS_AO112X4 U961 ( .A(n854), .B(n853), .C(n1018), .D(n852), .Z(n855) );
  HS65_GS_NAND2X2 U962 ( .A(n868), .B(n855), .Z(\mul_b2/result_sat[6] ) );
  HS65_GSS_XOR2X3 U963 ( .A(n857), .B(n856), .Z(n860) );
  HS65_GS_OAI21X2 U964 ( .A(n859), .B(n860), .C(n1034), .Z(n858) );
  HS65_GS_CBI4I1X3 U965 ( .A(n860), .B(n859), .C(n858), .D(n868), .Z(
        \mul_b2/result_sat[5] ) );
  HS65_GS_AOI12X2 U966 ( .A(n863), .B(n862), .C(n1033), .Z(n861) );
  HS65_GS_CBI4I6X2 U967 ( .A(n863), .B(n862), .C(n861), .D(n1018), .Z(
        \mul_b2/result_sat[1] ) );
  HS65_GS_AO112X4 U968 ( .A(n866), .B(n865), .C(n1018), .D(n864), .Z(n867) );
  HS65_GS_NAND2X2 U969 ( .A(n868), .B(n867), .Z(\mul_b2/result_sat[0] ) );
  HS65_GS_IVX2 U970 ( .A(n869), .Z(n871) );
  HS65_GS_AOI22X1 U971 ( .A(n872), .B(n871), .C(n873), .D(n870), .Z(n887) );
  HS65_GS_AOI12X2 U972 ( .A(n875), .B(n874), .C(n873), .Z(n885) );
  HS65_GS_FA1X4 U973 ( .A0(n878), .B0(n877), .CI(n876), .CO(n879), .S0(n884)
         );
  HS65_GS_FA1X4 U974 ( .A0(n881), .B0(n880), .CI(n879), .CO(n342), .S0(n883)
         );
  HS65_GS_NOR3X1 U975 ( .A(n885), .B(n884), .C(n883), .Z(n882) );
  HS65_GS_AOI12X2 U976 ( .A(n887), .B(n882), .C(\mul_b0/result_sat[15] ), .Z(
        n1056) );
  HS65_GS_IVX2 U977 ( .A(n1056), .Z(n939) );
  HS65_GS_NAND3X2 U978 ( .A(n885), .B(n884), .C(n883), .Z(n886) );
  HS65_GS_OAI21X2 U979 ( .A(n887), .B(n886), .C(\mul_b0/result_sat[15] ), .Z(
        n1053) );
  HS65_GS_IVX2 U980 ( .A(n1053), .Z(n1055) );
  HS65_GS_AO112X4 U981 ( .A(n890), .B(n889), .C(n1055), .D(n888), .Z(n891) );
  HS65_GS_NAND2X2 U982 ( .A(n939), .B(n891), .Z(\mul_b0/result_sat[12] ) );
  HS65_GS_AO112X4 U983 ( .A(n894), .B(n893), .C(n1055), .D(n892), .Z(n895) );
  HS65_GS_NAND2X2 U984 ( .A(n939), .B(n895), .Z(\mul_b0/result_sat[11] ) );
  HS65_GS_AO112X4 U985 ( .A(n898), .B(n897), .C(n1055), .D(n896), .Z(n899) );
  HS65_GS_NAND2X2 U986 ( .A(n939), .B(n899), .Z(\mul_b0/result_sat[10] ) );
  HS65_GS_AO112X4 U987 ( .A(n902), .B(n901), .C(n1055), .D(n900), .Z(n903) );
  HS65_GS_NAND2X2 U988 ( .A(n939), .B(n903), .Z(\mul_b0/result_sat[9] ) );
  HS65_GS_AO112X4 U989 ( .A(n906), .B(n905), .C(n1055), .D(n904), .Z(n907) );
  HS65_GS_NAND2X2 U990 ( .A(n939), .B(n907), .Z(\mul_b0/result_sat[8] ) );
  HS65_GS_AO112X4 U991 ( .A(n910), .B(n909), .C(n1055), .D(n908), .Z(n911) );
  HS65_GS_NAND2X2 U992 ( .A(n939), .B(n911), .Z(\mul_b0/result_sat[7] ) );
  HS65_GS_AO112X4 U993 ( .A(n914), .B(n913), .C(n1055), .D(n912), .Z(n915) );
  HS65_GS_NAND2X2 U994 ( .A(n939), .B(n915), .Z(\mul_b0/result_sat[6] ) );
  HS65_GS_AO112X4 U995 ( .A(n918), .B(n917), .C(n1055), .D(n916), .Z(n919) );
  HS65_GS_NAND2X2 U996 ( .A(n939), .B(n919), .Z(\mul_b0/result_sat[5] ) );
  HS65_GS_AO112X4 U997 ( .A(n922), .B(n921), .C(n1055), .D(n920), .Z(n923) );
  HS65_GS_NAND2X2 U998 ( .A(n939), .B(n923), .Z(\mul_b0/result_sat[4] ) );
  HS65_GS_AO112X4 U999 ( .A(n926), .B(n925), .C(n1055), .D(n924), .Z(n927) );
  HS65_GS_NAND2X2 U1000 ( .A(n939), .B(n927), .Z(\mul_b0/result_sat[3] ) );
  HS65_GS_AOI12X2 U1001 ( .A(n930), .B(n929), .C(n1056), .Z(n928) );
  HS65_GS_CBI4I6X2 U1002 ( .A(n930), .B(n929), .C(n928), .D(n1055), .Z(
        \mul_b0/result_sat[2] ) );
  HS65_GS_AO112X4 U1003 ( .A(n933), .B(n932), .C(n1055), .D(n931), .Z(n934) );
  HS65_GS_NAND2X2 U1004 ( .A(n939), .B(n934), .Z(\mul_b0/result_sat[1] ) );
  HS65_GS_AO112X4 U1005 ( .A(n937), .B(n936), .C(n1055), .D(n935), .Z(n938) );
  HS65_GS_NAND2X2 U1006 ( .A(n939), .B(n938), .Z(\mul_b0/result_sat[0] ) );
  HS65_GS_IVX2 U1007 ( .A(n1365), .Z(n1791) );
  HS65_GS_MUX21I1X3 U1008 ( .D0(n1661), .D1(data_out[2]), .S0(n1366), .Z(n1881) );
  HS65_GS_MUX21I1X3 U1009 ( .D0(n1659), .D1(data_out[3]), .S0(valid_in), .Z(
        n1878) );
  HS65_GS_MUX21I1X3 U1010 ( .D0(n1657), .D1(data_out[4]), .S0(n1792), .Z(n1875) );
  HS65_GS_MUX21I1X3 U1011 ( .D0(n1655), .D1(data_out[5]), .S0(n1366), .Z(n1872) );
  HS65_GS_MUX21I1X3 U1012 ( .D0(n1653), .D1(data_out[6]), .S0(valid_in), .Z(
        n1869) );
  HS65_GS_MUX21I1X3 U1013 ( .D0(n1651), .D1(data_out[7]), .S0(n1792), .Z(n1866) );
  HS65_GS_MUX21I1X3 U1014 ( .D0(n1649), .D1(data_out[8]), .S0(n1366), .Z(n1863) );
  HS65_GS_MUX21I1X3 U1015 ( .D0(n1647), .D1(data_out[9]), .S0(n1792), .Z(n1860) );
  HS65_GS_MUX21I1X3 U1016 ( .D0(n1645), .D1(data_out[10]), .S0(valid_in), .Z(
        n1857) );
  HS65_GS_MUX21I1X3 U1017 ( .D0(n1643), .D1(data_out[11]), .S0(n1366), .Z(
        n1854) );
  HS65_GS_MUX21I1X3 U1018 ( .D0(n1637), .D1(data_out[14]), .S0(n1792), .Z(
        n1845) );
  HS65_GS_MUX21I1X3 U1019 ( .D0(n1713), .D1(data_out[1]), .S0(n1792), .Z(n1884) );
  HS65_GS_MUX21I1X3 U1020 ( .D0(n1365), .D1(data_in[15]), .S0(n1792), .Z(n1793) );
  HS65_GS_IVX2 U1021 ( .A(n1710), .Z(n1790) );
  HS65_GS_BFX4 U1022 ( .A(n1792), .Z(n1382) );
  HS65_GS_MUX21I1X3 U1023 ( .D0(n1712), .D1(data_out[0]), .S0(n1382), .Z(n1887) );
  HS65_GSS_XNOR2X3 U1024 ( .A(n941), .B(n940), .Z(n963) );
  HS65_GS_IVX2 U1025 ( .A(n942), .Z(n962) );
  HS65_GS_FA1X4 U1026 ( .A0(n945), .B0(n944), .CI(n943), .CO(n947), .S0(n960)
         );
  HS65_GS_FA1X4 U1027 ( .A0(n948), .B0(n947), .CI(n946), .CO(n806), .S0(n958)
         );
  HS65_GS_FA1X4 U1028 ( .A0(n951), .B0(n950), .CI(n949), .CO(n953), .S0(n957)
         );
  HS65_GS_FA1X4 U1029 ( .A0(n954), .B0(n953), .CI(n952), .CO(n944), .S0(n956)
         );
  HS65_GS_OR3X4 U1030 ( .A(n958), .B(n957), .C(n956), .Z(n955) );
  HS65_GS_OAI21X2 U1031 ( .A(n960), .B(n955), .C(\mul_a1/result_sat[15] ), .Z(
        n1447) );
  HS65_GS_OAI21X2 U1032 ( .A(n962), .B(n963), .C(n1447), .Z(n961) );
  HS65_GS_AND3X4 U1033 ( .A(n958), .B(n957), .C(n956), .Z(n959) );
  HS65_GS_AOI12X2 U1034 ( .A(n960), .B(n959), .C(\mul_a1/result_sat[15] ), .Z(
        n1449) );
  HS65_GS_IVX2 U1035 ( .A(n1449), .Z(n1745) );
  HS65_GS_CBI4I1X3 U1036 ( .A(n963), .B(n962), .C(n961), .D(n1745), .Z(
        \mul_a1/result_sat[13] ) );
  HS65_GSS_XNOR2X3 U1037 ( .A(n965), .B(n964), .Z(n968) );
  HS65_GS_OAI21X2 U1038 ( .A(n967), .B(n968), .C(n1447), .Z(n966) );
  HS65_GS_CBI4I1X3 U1039 ( .A(n968), .B(n967), .C(n966), .D(n1745), .Z(
        \mul_a1/result_sat[8] ) );
  HS65_GS_OAI21X2 U1040 ( .A(n970), .B(n971), .C(n1447), .Z(n969) );
  HS65_GS_CBI4I1X3 U1041 ( .A(n971), .B(n970), .C(n969), .D(n1745), .Z(
        \mul_a1/result_sat[7] ) );
  HS65_GS_OAI21X2 U1042 ( .A(n973), .B(n974), .C(n1447), .Z(n972) );
  HS65_GS_CBI4I1X3 U1043 ( .A(n974), .B(n973), .C(n972), .D(n1745), .Z(
        \mul_a1/result_sat[5] ) );
  HS65_GS_OAI21X2 U1044 ( .A(n976), .B(n977), .C(n1447), .Z(n975) );
  HS65_GS_CBI4I1X3 U1045 ( .A(n977), .B(n976), .C(n975), .D(n1745), .Z(
        \mul_a1/result_sat[4] ) );
  HS65_GS_OAI21X2 U1046 ( .A(n979), .B(n980), .C(n1447), .Z(n978) );
  HS65_GS_CBI4I1X3 U1047 ( .A(n980), .B(n979), .C(n978), .D(n1745), .Z(
        \mul_a1/result_sat[2] ) );
  HS65_GS_NOR2X2 U1048 ( .A(n1726), .B(n1727), .Z(\mul_b2/fa1_c0[17] ) );
  HS65_GS_NOR2X2 U1049 ( .A(n1725), .B(n1728), .Z(\mul_b2/fa1_c0[16] ) );
  HS65_GS_NOR2X2 U1050 ( .A(n1724), .B(n1726), .Z(\mul_b2/fa1_c0[15] ) );
  HS65_GS_NOR2X2 U1051 ( .A(n1723), .B(n1725), .Z(\mul_b2/fa1_c0[14] ) );
  HS65_GS_NOR2X2 U1052 ( .A(n1722), .B(n1724), .Z(\mul_b2/fa1_c0[13] ) );
  HS65_GS_NOR2X2 U1053 ( .A(n1721), .B(n1723), .Z(\mul_b2/fa1_c0[12] ) );
  HS65_GS_NOR2X2 U1054 ( .A(n1720), .B(n1722), .Z(\mul_b2/fa1_c0[11] ) );
  HS65_GS_NOR2X2 U1055 ( .A(n1719), .B(n1721), .Z(\mul_b2/fa1_c0[10] ) );
  HS65_GS_NOR2X2 U1056 ( .A(n1718), .B(n1720), .Z(\mul_b2/fa1_c0[9] ) );
  HS65_GS_NOR2X2 U1057 ( .A(n1717), .B(n1719), .Z(\mul_b2/fa1_c0[8] ) );
  HS65_GS_NOR2X2 U1058 ( .A(n1716), .B(n1718), .Z(\mul_b2/fa1_c0[7] ) );
  HS65_GS_NOR2X2 U1059 ( .A(n1715), .B(n1717), .Z(\mul_b2/fa1_c0[6] ) );
  HS65_GS_NOR2X2 U1060 ( .A(n1714), .B(n1716), .Z(\mul_b2/fa1_c0[5] ) );
  HS65_GS_IVX2 U1061 ( .A(n1727), .Z(n1789) );
  HS65_GS_IVX2 U1062 ( .A(y_z2[14]), .Z(n1510) );
  HS65_GS_IVX2 U1063 ( .A(y_z2[13]), .Z(n1512) );
  HS65_GS_IVX2 U1064 ( .A(y_z2[12]), .Z(n1514) );
  HS65_GS_IVX2 U1065 ( .A(y_z2[11]), .Z(n1516) );
  HS65_GS_IVX2 U1066 ( .A(y_z2[10]), .Z(n1518) );
  HS65_GS_IVX2 U1067 ( .A(y_z2[9]), .Z(n1520) );
  HS65_GS_IVX2 U1068 ( .A(y_z2[8]), .Z(n1522) );
  HS65_GS_IVX2 U1069 ( .A(y_z2[7]), .Z(n1524) );
  HS65_GS_IVX2 U1070 ( .A(y_z2[6]), .Z(n1526) );
  HS65_GS_IVX2 U1071 ( .A(y_z2[5]), .Z(n1528) );
  HS65_GS_IVX2 U1072 ( .A(y_z2[4]), .Z(n1530) );
  HS65_GS_IVX2 U1073 ( .A(y_z2[3]), .Z(n1532) );
  HS65_GS_IVX2 U1074 ( .A(y_z2[2]), .Z(n1534) );
  HS65_GS_IVX2 U1075 ( .A(y_z2[1]), .Z(n1708) );
  HS65_GS_IVX2 U1076 ( .A(y_z2[0]), .Z(n1707) );
  HS65_GS_NOR2X2 U1077 ( .A(y_z2[15]), .B(n1455), .Z(n1785) );
  HS65_GSS_XOR2X3 U1078 ( .A(n1785), .B(n981), .Z(\mul_a2/fa1_s1[23] ) );
  HS65_GS_NOR2X2 U1079 ( .A(n1728), .B(n1727), .Z(\mul_b2/fa1_c0[18] ) );
  HS65_GS_NOR2X2 U1080 ( .A(x_z2[15]), .B(n990), .Z(n982) );
  HS65_GSS_XNOR2X3 U1081 ( .A(n982), .B(n1680), .Z(\mul_b1/fa1_s1[27] ) );
  HS65_GS_IVX2 U1082 ( .A(x_z2[1]), .Z(n1349) );
  HS65_GS_IVX2 U1083 ( .A(x_z2[0]), .Z(n1347) );
  HS65_GS_NOR2X2 U1084 ( .A(x_z2[15]), .B(n1036), .Z(n983) );
  HS65_GSS_XNOR2X3 U1085 ( .A(n983), .B(n1680), .Z(\mul_b1/fa1_s2[29] ) );
  HS65_GS_IVX2 U1086 ( .A(x_z1[14]), .Z(n1364) );
  HS65_GS_IVX2 U1087 ( .A(x_z1[13]), .Z(n1363) );
  HS65_GS_IVX2 U1088 ( .A(x_z1[12]), .Z(n1362) );
  HS65_GS_IVX2 U1089 ( .A(x_z1[11]), .Z(n1360) );
  HS65_GS_IVX2 U1090 ( .A(x_z1[10]), .Z(n1359) );
  HS65_GS_IVX2 U1091 ( .A(x_z1[9]), .Z(n1358) );
  HS65_GS_IVX2 U1092 ( .A(x_z1[8]), .Z(n1357) );
  HS65_GS_IVX2 U1093 ( .A(x_z1[7]), .Z(n1356) );
  HS65_GS_IVX2 U1094 ( .A(x_z1[6]), .Z(n1355) );
  HS65_GS_IVX2 U1095 ( .A(x_z1[5]), .Z(n1354) );
  HS65_GS_IVX2 U1096 ( .A(x_z1[4]), .Z(n1353) );
  HS65_GS_IVX2 U1097 ( .A(x_z1[3]), .Z(n1352) );
  HS65_GS_IVX2 U1098 ( .A(x_z1[2]), .Z(n1351) );
  HS65_GS_IVX2 U1099 ( .A(x_z1[1]), .Z(n1350) );
  HS65_GS_IVX2 U1100 ( .A(x_z1[0]), .Z(n1348) );
  HS65_GS_NOR2X2 U1101 ( .A(n1791), .B(n985), .Z(n984) );
  HS65_GSS_XNOR2X3 U1102 ( .A(n984), .B(n1365), .Z(\mul_b0/fa1_s0[31] ) );
  HS65_GSS_XNOR2X3 U1103 ( .A(x_z1[15]), .B(n985), .Z(n1145) );
  HS65_GSS_XNOR2X3 U1104 ( .A(n1145), .B(n1365), .Z(\mul_b0/fa1_s0[20] ) );
  HS65_GS_NOR2X2 U1105 ( .A(y_z1[15]), .B(n1402), .Z(n1416) );
  HS65_GSS_XNOR2X3 U1106 ( .A(n1416), .B(n1635), .Z(\mul_a1/fa1_s1[29] ) );
  HS65_GSS_XNOR2X3 U1107 ( .A(n1416), .B(n1637), .Z(\mul_a1/fa1_s1[25] ) );
  HS65_GS_NOR2X2 U1108 ( .A(n1790), .B(n1367), .Z(n986) );
  HS65_GSS_XNOR2X3 U1109 ( .A(n986), .B(n1710), .Z(\mul_a2/fa1_s2[29] ) );
  HS65_GSS_XNOR2X3 U1110 ( .A(n1632), .B(n1637), .Z(\mul_a1/fa1_s0[17] ) );
  HS65_GS_HA1X4 U1111 ( .A0(n1682), .B0(n987), .CO(n991), .S0(n992) );
  HS65_GS_AND2X4 U1112 ( .A(n992), .B(x_z2[12]), .Z(\mul_b1/fa1_c1[20] ) );
  HS65_GS_HA1X4 U1113 ( .A0(n1692), .B0(n988), .CO(n989), .S0(n997) );
  HS65_GS_AND2X4 U1114 ( .A(n997), .B(x_z2[7]), .Z(\mul_b1/fa1_c1[15] ) );
  HS65_GS_HA1X4 U1115 ( .A0(n1690), .B0(n989), .CO(n995), .S0(n996) );
  HS65_GS_AND2X4 U1116 ( .A(n996), .B(x_z2[8]), .Z(\mul_b1/fa1_c1[16] ) );
  HS65_GSS_XNOR2X3 U1117 ( .A(x_z2[15]), .B(n990), .Z(n1007) );
  HS65_GSS_XNOR2X3 U1118 ( .A(n1007), .B(n1682), .Z(\mul_b1/fa1_s1[22] ) );
  HS65_GS_HA1X4 U1119 ( .A0(n1680), .B0(n991), .CO(n990), .S0(n1008) );
  HS65_GSS_XNOR2X3 U1120 ( .A(n1008), .B(n1684), .Z(\mul_b1/fa1_s1[21] ) );
  HS65_GSS_XNOR2X3 U1121 ( .A(n992), .B(n1686), .Z(\mul_b1/fa1_s1[20] ) );
  HS65_GS_HA1X4 U1122 ( .A0(n1684), .B0(n993), .CO(n987), .S0(n1009) );
  HS65_GSS_XNOR2X3 U1123 ( .A(n1009), .B(n1688), .Z(\mul_b1/fa1_s1[19] ) );
  HS65_GS_HA1X4 U1124 ( .A0(n1686), .B0(n994), .CO(n993), .S0(n1006) );
  HS65_GSS_XNOR2X3 U1125 ( .A(n1006), .B(n1690), .Z(\mul_b1/fa1_s1[18] ) );
  HS65_GS_HA1X4 U1126 ( .A0(n1688), .B0(n995), .CO(n994), .S0(n1004) );
  HS65_GSS_XNOR2X3 U1127 ( .A(n1004), .B(n1692), .Z(\mul_b1/fa1_s1[17] ) );
  HS65_GSS_XNOR2X3 U1128 ( .A(n996), .B(n1694), .Z(\mul_b1/fa1_s1[16] ) );
  HS65_GSS_XNOR2X3 U1129 ( .A(n997), .B(n1696), .Z(\mul_b1/fa1_s1[15] ) );
  HS65_GS_HA1X4 U1130 ( .A0(n1694), .B0(n998), .CO(n988), .S0(n1131) );
  HS65_GSS_XNOR2X3 U1131 ( .A(n1131), .B(n1698), .Z(\mul_b1/fa1_s1[14] ) );
  HS65_GS_HA1X4 U1132 ( .A0(n1696), .B0(n999), .CO(n998), .S0(n1060) );
  HS65_GSS_XNOR2X3 U1133 ( .A(n1060), .B(n1700), .Z(\mul_b1/fa1_s1[13] ) );
  HS65_GS_HA1X4 U1134 ( .A0(n1698), .B0(n1000), .CO(n999), .S0(n1061) );
  HS65_GSS_XNOR2X3 U1135 ( .A(n1061), .B(n1702), .Z(\mul_b1/fa1_s1[12] ) );
  HS65_GS_HA1X4 U1136 ( .A0(n1700), .B0(n1001), .CO(n1000), .S0(n1062) );
  HS65_GSS_XNOR2X3 U1137 ( .A(n1062), .B(n1704), .Z(\mul_b1/fa1_s1[11] ) );
  HS65_GS_HA1X4 U1138 ( .A0(n1702), .B0(n1002), .CO(n1001), .S0(n1063) );
  HS65_GSS_XNOR2X3 U1139 ( .A(n1063), .B(n1706), .Z(\mul_b1/fa1_s1[10] ) );
  HS65_GS_HA1X4 U1140 ( .A0(n1704), .B0(n1003), .CO(n1002), .S0(n1064) );
  HS65_GSS_XNOR2X3 U1141 ( .A(n1064), .B(n1349), .Z(\mul_b1/fa1_s1[9] ) );
  HS65_GS_AND2X4 U1142 ( .A(n1004), .B(x_z2[9]), .Z(\mul_b1/fa1_c1[17] ) );
  HS65_GS_HA1X4 U1143 ( .A0(n1706), .B0(n1005), .CO(n1003), .S0(n1065) );
  HS65_GSS_XNOR2X3 U1144 ( .A(n1065), .B(n1347), .Z(\mul_b1/fa1_s1[8] ) );
  HS65_GS_AND2X4 U1145 ( .A(n1006), .B(x_z2[10]), .Z(\mul_b1/fa1_c1[18] ) );
  HS65_GS_AND2X4 U1146 ( .A(n1007), .B(x_z2[14]), .Z(\mul_b1/fa1_c1[22] ) );
  HS65_GS_AND2X4 U1147 ( .A(n1008), .B(x_z2[13]), .Z(\mul_b1/fa1_c1[21] ) );
  HS65_GS_AND2X4 U1148 ( .A(n1009), .B(x_z2[11]), .Z(\mul_b1/fa1_c1[19] ) );
  HS65_GS_FA1X4 U1149 ( .A0(n1012), .B0(n1011), .CI(n1010), .CO(n819), .S0(
        n1013) );
  HS65_GS_AO12X4 U1150 ( .A(n1013), .B(n1034), .C(n1033), .Z(
        \mul_b2/result_sat[14] ) );
  HS65_GS_FA1X4 U1151 ( .A0(n1016), .B0(n1015), .CI(n1014), .CO(n1010), .S0(
        n1017) );
  HS65_GS_OA12X4 U1152 ( .A(n1033), .B(n1017), .C(n1034), .Z(
        \mul_b2/result_sat[13] ) );
  HS65_GS_AOI12X2 U1153 ( .A(n1021), .B(n1020), .C(n1018), .Z(n1019) );
  HS65_GS_CB4I6X4 U1154 ( .A(n1021), .B(n1020), .C(n1019), .D(n1033), .Z(
        \mul_b2/result_sat[12] ) );
  HS65_GS_FA1X4 U1155 ( .A0(n1024), .B0(n1023), .CI(n1022), .CO(n859), .S0(
        n1025) );
  HS65_GS_OA12X4 U1156 ( .A(n1033), .B(n1025), .C(n1034), .Z(
        \mul_b2/result_sat[4] ) );
  HS65_GS_FA1X4 U1157 ( .A0(n1028), .B0(n1027), .CI(n1026), .CO(n1024), .S0(
        n1029) );
  HS65_GS_AO12X4 U1158 ( .A(n1029), .B(n1034), .C(n1033), .Z(
        \mul_b2/result_sat[3] ) );
  HS65_GS_FA1X4 U1159 ( .A0(n1032), .B0(n1031), .CI(n1030), .CO(n1026), .S0(
        n1035) );
  HS65_GS_AO12X4 U1160 ( .A(n1035), .B(n1034), .C(n1033), .Z(
        \mul_b2/result_sat[2] ) );
  HS65_GSS_XNOR2X3 U1161 ( .A(x_z2[15]), .B(n1036), .Z(n1066) );
  HS65_GS_AND2X4 U1162 ( .A(n1066), .B(x_z2[14]), .Z(\mul_b1/fa1_c2[28] ) );
  HS65_GS_HA1X4 U1163 ( .A0(n1682), .B0(n1037), .CO(n1036), .S0(n1067) );
  HS65_GS_AND2X4 U1164 ( .A(n1067), .B(x_z2[13]), .Z(\mul_b1/fa1_c2[27] ) );
  HS65_GS_HA1X4 U1165 ( .A0(n1684), .B0(n1038), .CO(n1037), .S0(n1068) );
  HS65_GS_AND2X4 U1166 ( .A(n1068), .B(x_z2[12]), .Z(\mul_b1/fa1_c2[26] ) );
  HS65_GS_HA1X4 U1167 ( .A0(n1686), .B0(n1039), .CO(n1038), .S0(n1069) );
  HS65_GS_AND2X4 U1168 ( .A(n1069), .B(x_z2[11]), .Z(\mul_b1/fa1_c2[25] ) );
  HS65_GS_HA1X4 U1169 ( .A0(n1688), .B0(n1040), .CO(n1039), .S0(n1070) );
  HS65_GS_AND2X4 U1170 ( .A(n1070), .B(x_z2[10]), .Z(\mul_b1/fa1_c2[24] ) );
  HS65_GS_HA1X4 U1171 ( .A0(n1690), .B0(n1041), .CO(n1040), .S0(n1071) );
  HS65_GS_AND2X4 U1172 ( .A(n1071), .B(x_z2[9]), .Z(\mul_b1/fa1_c2[23] ) );
  HS65_GS_HA1X4 U1173 ( .A0(n1692), .B0(n1042), .CO(n1041), .S0(n1072) );
  HS65_GS_AND2X4 U1174 ( .A(n1072), .B(x_z2[8]), .Z(\mul_b1/fa1_c2[22] ) );
  HS65_GS_HA1X4 U1175 ( .A0(n1694), .B0(n1043), .CO(n1042), .S0(n1073) );
  HS65_GS_AND2X4 U1176 ( .A(n1073), .B(x_z2[7]), .Z(\mul_b1/fa1_c2[21] ) );
  HS65_GS_HA1X4 U1177 ( .A0(n1696), .B0(n1044), .CO(n1043), .S0(n1074) );
  HS65_GS_AND2X4 U1178 ( .A(n1074), .B(x_z2[6]), .Z(\mul_b1/fa1_c2[20] ) );
  HS65_GS_HA1X4 U1179 ( .A0(n1698), .B0(n1045), .CO(n1044), .S0(n1075) );
  HS65_GS_AND2X4 U1180 ( .A(n1075), .B(x_z2[5]), .Z(\mul_b1/fa1_c2[19] ) );
  HS65_GS_HA1X4 U1181 ( .A0(n1700), .B0(n1046), .CO(n1045), .S0(n1076) );
  HS65_GS_AND2X4 U1182 ( .A(n1076), .B(x_z2[4]), .Z(\mul_b1/fa1_c2[18] ) );
  HS65_GS_HA1X4 U1183 ( .A0(n1702), .B0(n1047), .CO(n1046), .S0(n1077) );
  HS65_GS_AND2X4 U1184 ( .A(n1077), .B(x_z2[3]), .Z(\mul_b1/fa1_c2[17] ) );
  HS65_GS_HA1X4 U1185 ( .A0(n1704), .B0(n1048), .CO(n1047), .S0(n1078) );
  HS65_GS_AND2X4 U1186 ( .A(n1078), .B(x_z2[2]), .Z(\mul_b1/fa1_c2[16] ) );
  HS65_GS_HA1X4 U1187 ( .A0(n1706), .B0(n1049), .CO(n1048), .S0(n1079) );
  HS65_GS_AND2X4 U1188 ( .A(n1079), .B(x_z2[1]), .Z(\mul_b1/fa1_c2[15] ) );
  HS65_GS_HA1X4 U1189 ( .A0(n1349), .B0(n1347), .CO(n1049), .S0(n1080) );
  HS65_GS_AND2X4 U1190 ( .A(n1080), .B(x_z2[0]), .Z(\mul_b1/fa1_c2[14] ) );
  HS65_GS_FA1X4 U1191 ( .A0(n1052), .B0(n1051), .CI(n1050), .CO(n876), .S0(
        n1054) );
  HS65_GS_AO12X4 U1192 ( .A(n1054), .B(n1053), .C(n1056), .Z(
        \mul_b0/result_sat[14] ) );
  HS65_GS_AOI12X2 U1193 ( .A(n1059), .B(n1058), .C(n1055), .Z(n1057) );
  HS65_GS_CB4I6X4 U1194 ( .A(n1059), .B(n1058), .C(n1057), .D(n1056), .Z(
        \mul_b0/result_sat[13] ) );
  HS65_GS_AND2X4 U1195 ( .A(n1060), .B(x_z2[5]), .Z(\mul_b1/fa1_c1[13] ) );
  HS65_GS_AND2X4 U1196 ( .A(n1061), .B(x_z2[4]), .Z(\mul_b1/fa1_c1[12] ) );
  HS65_GS_AND2X4 U1197 ( .A(n1062), .B(x_z2[3]), .Z(\mul_b1/fa1_c1[11] ) );
  HS65_GS_AND2X4 U1198 ( .A(n1063), .B(x_z2[2]), .Z(\mul_b1/fa1_c1[10] ) );
  HS65_GS_AND2X4 U1199 ( .A(n1064), .B(x_z2[1]), .Z(\mul_b1/fa1_c1[9] ) );
  HS65_GS_AND2X4 U1200 ( .A(n1065), .B(x_z2[0]), .Z(\mul_b1/fa1_c1[8] ) );
  HS65_GSS_XNOR2X3 U1201 ( .A(n1066), .B(n1682), .Z(\mul_b1/fa1_s2[28] ) );
  HS65_GSS_XNOR2X3 U1202 ( .A(n1067), .B(n1684), .Z(\mul_b1/fa1_s2[27] ) );
  HS65_GSS_XNOR2X3 U1203 ( .A(n1068), .B(n1686), .Z(\mul_b1/fa1_s2[26] ) );
  HS65_GSS_XNOR2X3 U1204 ( .A(n1069), .B(n1688), .Z(\mul_b1/fa1_s2[25] ) );
  HS65_GSS_XNOR2X3 U1205 ( .A(n1070), .B(n1690), .Z(\mul_b1/fa1_s2[24] ) );
  HS65_GSS_XNOR2X3 U1206 ( .A(n1071), .B(n1692), .Z(\mul_b1/fa1_s2[23] ) );
  HS65_GSS_XNOR2X3 U1207 ( .A(n1072), .B(n1694), .Z(\mul_b1/fa1_s2[22] ) );
  HS65_GSS_XNOR2X3 U1208 ( .A(n1073), .B(n1696), .Z(\mul_b1/fa1_s2[21] ) );
  HS65_GSS_XNOR2X3 U1209 ( .A(n1074), .B(n1698), .Z(\mul_b1/fa1_s2[20] ) );
  HS65_GSS_XNOR2X3 U1210 ( .A(n1075), .B(n1700), .Z(\mul_b1/fa1_s2[19] ) );
  HS65_GSS_XNOR2X3 U1211 ( .A(n1076), .B(n1702), .Z(\mul_b1/fa1_s2[18] ) );
  HS65_GSS_XNOR2X3 U1212 ( .A(n1077), .B(n1704), .Z(\mul_b1/fa1_s2[17] ) );
  HS65_GSS_XNOR2X3 U1213 ( .A(n1078), .B(n1706), .Z(\mul_b1/fa1_s2[16] ) );
  HS65_GSS_XNOR2X3 U1214 ( .A(n1079), .B(n1349), .Z(\mul_b1/fa1_s2[15] ) );
  HS65_GSS_XNOR2X3 U1215 ( .A(n1080), .B(n1347), .Z(\mul_b1/fa1_s2[14] ) );
  HS65_GS_FA1X4 U1216 ( .A0(n1083), .B0(n1082), .CI(n1081), .CO(n1086), .S0(
        n1084) );
  HS65_GS_IVX2 U1217 ( .A(n1084), .Z(n1102) );
  HS65_GS_FA1X4 U1218 ( .A0(n1087), .B0(n1086), .CI(n1085), .CO(n1090), .S0(
        n1100) );
  HS65_GS_FA1X4 U1219 ( .A0(n1090), .B0(n1089), .CI(n1088), .CO(n533), .S0(
        n1099) );
  HS65_GS_FA1X4 U1220 ( .A0(n1093), .B0(n1092), .CI(n1091), .CO(n1083), .S0(
        n1098) );
  HS65_GS_NOR3X1 U1221 ( .A(n1100), .B(n1099), .C(n1098), .Z(n1094) );
  HS65_GS_AOI12X2 U1222 ( .A(n1102), .B(n1094), .C(\mul_b1/result_sat[15] ), 
        .Z(n1122) );
  HS65_GS_FA1X4 U1223 ( .A0(n1097), .B0(n1096), .CI(n1095), .CO(n1092), .S0(
        n1103) );
  HS65_GS_NAND3X2 U1224 ( .A(n1100), .B(n1099), .C(n1098), .Z(n1101) );
  HS65_GS_OAI21X2 U1225 ( .A(n1102), .B(n1101), .C(\mul_b1/result_sat[15] ), 
        .Z(n1750) );
  HS65_GS_OA12X4 U1226 ( .A(n1122), .B(n1103), .C(n1750), .Z(
        \mul_b1/result_sat[14] ) );
  HS65_GS_FA1X4 U1227 ( .A0(n1106), .B0(n1105), .CI(n1104), .CO(n1096), .S0(
        n1107) );
  HS65_GS_OA12X4 U1228 ( .A(n1122), .B(n1107), .C(n1750), .Z(
        \mul_b1/result_sat[13] ) );
  HS65_GS_FA1X4 U1229 ( .A0(n1110), .B0(n1109), .CI(n1108), .CO(n1106), .S0(
        n1111) );
  HS65_GS_OA12X4 U1230 ( .A(n1122), .B(n1111), .C(n1750), .Z(
        \mul_b1/result_sat[12] ) );
  HS65_GS_FA1X4 U1231 ( .A0(n1114), .B0(n1113), .CI(n1112), .CO(n1109), .S0(
        n1115) );
  HS65_GS_AO12X4 U1232 ( .A(n1115), .B(n1750), .C(n1122), .Z(
        \mul_b1/result_sat[11] ) );
  HS65_GS_FA1X4 U1233 ( .A0(n1118), .B0(n1117), .CI(n1116), .CO(n1113), .S0(
        n1119) );
  HS65_GS_AO12X4 U1234 ( .A(n1119), .B(n1750), .C(n1122), .Z(
        \mul_b1/result_sat[10] ) );
  HS65_GSS_XNOR2X3 U1235 ( .A(n1121), .B(n1120), .Z(n1124) );
  HS65_GS_IVX2 U1236 ( .A(n1122), .Z(n1780) );
  HS65_GS_OAI21X2 U1237 ( .A(n1124), .B(n1125), .C(n1780), .Z(n1123) );
  HS65_GS_CB4I1X4 U1238 ( .A(n1125), .B(n1124), .C(n1123), .D(n1750), .Z(
        \mul_b1/result_sat[9] ) );
  HS65_GSS_XNOR2X3 U1239 ( .A(n1127), .B(n1126), .Z(n1129) );
  HS65_GS_OAI21X2 U1240 ( .A(n1129), .B(n1130), .C(n1780), .Z(n1128) );
  HS65_GS_CB4I1X4 U1241 ( .A(n1130), .B(n1129), .C(n1128), .D(n1750), .Z(
        \mul_b1/result_sat[8] ) );
  HS65_GS_AND2X4 U1242 ( .A(n1131), .B(x_z2[6]), .Z(\mul_b1/fa1_c1[14] ) );
  HS65_GS_HA1X4 U1243 ( .A0(n1364), .B0(n1132), .CO(n985), .S0(n1146) );
  HS65_GSS_XNOR2X3 U1244 ( .A(n1146), .B(n1365), .Z(\mul_b0/fa1_s0[19] ) );
  HS65_GS_HA1X4 U1245 ( .A0(n1363), .B0(n1133), .CO(n1132), .S0(n1147) );
  HS65_GSS_XNOR2X3 U1246 ( .A(n1147), .B(n1365), .Z(\mul_b0/fa1_s0[18] ) );
  HS65_GS_HA1X4 U1247 ( .A0(n1362), .B0(n1134), .CO(n1133), .S0(n1148) );
  HS65_GSS_XNOR2X3 U1248 ( .A(n1148), .B(n1365), .Z(\mul_b0/fa1_s0[17] ) );
  HS65_GS_HA1X4 U1249 ( .A0(n1360), .B0(n1135), .CO(n1134), .S0(n1149) );
  HS65_GSS_XNOR2X3 U1250 ( .A(n1149), .B(n1365), .Z(\mul_b0/fa1_s0[16] ) );
  HS65_GS_HA1X4 U1251 ( .A0(n1359), .B0(n1136), .CO(n1135), .S0(n1150) );
  HS65_GSS_XNOR2X3 U1252 ( .A(n1150), .B(n1365), .Z(\mul_b0/fa1_s0[15] ) );
  HS65_GS_HA1X4 U1253 ( .A0(n1358), .B0(n1137), .CO(n1136), .S0(n1151) );
  HS65_GSS_XNOR2X3 U1254 ( .A(n1151), .B(n1364), .Z(\mul_b0/fa1_s0[14] ) );
  HS65_GS_HA1X4 U1255 ( .A0(n1357), .B0(n1138), .CO(n1137), .S0(n1152) );
  HS65_GSS_XNOR2X3 U1256 ( .A(n1152), .B(n1363), .Z(\mul_b0/fa1_s0[13] ) );
  HS65_GS_HA1X4 U1257 ( .A0(n1356), .B0(n1139), .CO(n1138), .S0(n1153) );
  HS65_GSS_XNOR2X3 U1258 ( .A(n1153), .B(n1362), .Z(\mul_b0/fa1_s0[12] ) );
  HS65_GS_HA1X4 U1259 ( .A0(n1355), .B0(n1140), .CO(n1139), .S0(n1154) );
  HS65_GSS_XNOR2X3 U1260 ( .A(n1154), .B(n1360), .Z(\mul_b0/fa1_s0[11] ) );
  HS65_GS_HA1X4 U1261 ( .A0(n1354), .B0(n1141), .CO(n1140), .S0(n1155) );
  HS65_GSS_XNOR2X3 U1262 ( .A(n1155), .B(n1359), .Z(\mul_b0/fa1_s0[10] ) );
  HS65_GS_HA1X4 U1263 ( .A0(n1353), .B0(n1142), .CO(n1141), .S0(n1156) );
  HS65_GSS_XNOR2X3 U1264 ( .A(n1156), .B(n1358), .Z(\mul_b0/fa1_s0[9] ) );
  HS65_GS_HA1X4 U1265 ( .A0(n1352), .B0(n1143), .CO(n1142), .S0(n1157) );
  HS65_GSS_XNOR2X3 U1266 ( .A(n1157), .B(n1357), .Z(\mul_b0/fa1_s0[8] ) );
  HS65_GS_HA1X4 U1267 ( .A0(n1351), .B0(n1144), .CO(n1143), .S0(n1158) );
  HS65_GSS_XNOR2X3 U1268 ( .A(n1158), .B(n1356), .Z(\mul_b0/fa1_s0[7] ) );
  HS65_GS_HA1X4 U1269 ( .A0(n1350), .B0(n1348), .CO(n1144), .S0(n1159) );
  HS65_GSS_XNOR2X3 U1270 ( .A(n1159), .B(n1355), .Z(\mul_b0/fa1_s0[6] ) );
  HS65_GS_AND2X4 U1271 ( .A(n1145), .B(n1791), .Z(\mul_b0/fa1_c0[20] ) );
  HS65_GS_AND2X4 U1272 ( .A(n1146), .B(x_z1[15]), .Z(\mul_b0/fa1_c0[19] ) );
  HS65_GS_AND2X4 U1273 ( .A(n1147), .B(n1791), .Z(\mul_b0/fa1_c0[18] ) );
  HS65_GS_AND2X4 U1274 ( .A(n1148), .B(x_z1[15]), .Z(\mul_b0/fa1_c0[17] ) );
  HS65_GS_AND2X4 U1275 ( .A(n1149), .B(n1791), .Z(\mul_b0/fa1_c0[16] ) );
  HS65_GS_AND2X4 U1276 ( .A(n1150), .B(x_z1[15]), .Z(\mul_b0/fa1_c0[15] ) );
  HS65_GS_AND2X4 U1277 ( .A(n1151), .B(x_z1[14]), .Z(\mul_b0/fa1_c0[14] ) );
  HS65_GS_AND2X4 U1278 ( .A(n1152), .B(x_z1[13]), .Z(\mul_b0/fa1_c0[13] ) );
  HS65_GS_AND2X4 U1279 ( .A(n1153), .B(x_z1[12]), .Z(\mul_b0/fa1_c0[12] ) );
  HS65_GS_AND2X4 U1280 ( .A(n1154), .B(x_z1[11]), .Z(\mul_b0/fa1_c0[11] ) );
  HS65_GS_AND2X4 U1281 ( .A(n1155), .B(x_z1[10]), .Z(\mul_b0/fa1_c0[10] ) );
  HS65_GS_AND2X4 U1282 ( .A(n1156), .B(x_z1[9]), .Z(\mul_b0/fa1_c0[9] ) );
  HS65_GS_AND2X4 U1283 ( .A(n1157), .B(x_z1[8]), .Z(\mul_b0/fa1_c0[8] ) );
  HS65_GS_AND2X4 U1284 ( .A(n1158), .B(x_z1[7]), .Z(\mul_b0/fa1_c0[7] ) );
  HS65_GS_AND2X4 U1285 ( .A(x_z1[6]), .B(n1159), .Z(\mul_b0/fa1_c0[6] ) );
  HS65_GS_AND2X4 U1286 ( .A(x_z1[5]), .B(x_z1[0]), .Z(\mul_b0/fa1_c0[5] ) );
  HS65_GS_IVX2 U1287 ( .A(valid_T3), .Z(n1784) );
  HS65_GS_AND2X4 U1288 ( .A(p_b1[1]), .B(p_b0[1]), .Z(n1203) );
  HS65_GSS_XOR2X3 U1289 ( .A(p_b1[1]), .B(p_b0[1]), .Z(n1206) );
  HS65_GS_FA1X4 U1290 ( .A0(p_b0[2]), .B0(p_b1[2]), .CI(p_b2[2]), .CO(n1199), 
        .S0(n1201) );
  HS65_GS_FA1X4 U1291 ( .A0(p_b0[3]), .B0(p_b1[3]), .CI(p_b2[3]), .CO(n1195), 
        .S0(n1197) );
  HS65_GS_FA1X4 U1292 ( .A0(p_b0[4]), .B0(p_b1[4]), .CI(p_b2[4]), .CO(n1191), 
        .S0(n1193) );
  HS65_GS_FA1X4 U1293 ( .A0(p_b0[5]), .B0(p_b1[5]), .CI(p_b2[5]), .CO(n1187), 
        .S0(n1189) );
  HS65_GS_FA1X4 U1294 ( .A0(p_b0[6]), .B0(p_b1[6]), .CI(p_b2[6]), .CO(n1183), 
        .S0(n1185) );
  HS65_GS_FA1X4 U1295 ( .A0(p_b0[7]), .B0(p_b1[7]), .CI(p_b2[7]), .CO(n1179), 
        .S0(n1181) );
  HS65_GS_FA1X4 U1296 ( .A0(p_b0[8]), .B0(p_b1[8]), .CI(p_b2[8]), .CO(n1175), 
        .S0(n1177) );
  HS65_GS_FA1X4 U1297 ( .A0(p_b0[9]), .B0(p_b1[9]), .CI(p_b2[9]), .CO(n1171), 
        .S0(n1173) );
  HS65_GS_FA1X4 U1298 ( .A0(p_b0[10]), .B0(p_b1[10]), .CI(p_b2[10]), .CO(n1163), .S0(n1169) );
  HS65_GS_FA1X4 U1299 ( .A0(p_b0[11]), .B0(p_b1[11]), .CI(p_b2[11]), .CO(n1167), .S0(n1161) );
  HS65_GS_FA1X4 U1300 ( .A0(p_b0[12]), .B0(p_b1[12]), .CI(p_b2[12]), .CO(n1256), .S0(n1165) );
  HS65_GS_IVX2 U1301 ( .A(n1160), .Z(n1253) );
  HS65_GS_FA1X4 U1302 ( .A0(n1163), .B0(n1162), .CI(n1161), .CO(n1166), .S0(
        n1164) );
  HS65_GS_IVX2 U1303 ( .A(n1164), .Z(n1246) );
  HS65_GS_FA1X4 U1304 ( .A0(n1167), .B0(n1166), .CI(n1165), .CO(n1255), .S0(
        n1168) );
  HS65_GS_IVX2 U1305 ( .A(n1168), .Z(n1250) );
  HS65_GS_FA1X4 U1306 ( .A0(n1171), .B0(n1170), .CI(n1169), .CO(n1162), .S0(
        n1172) );
  HS65_GS_IVX2 U1307 ( .A(n1172), .Z(n1242) );
  HS65_GS_FA1X4 U1308 ( .A0(n1175), .B0(n1174), .CI(n1173), .CO(n1170), .S0(
        n1176) );
  HS65_GS_IVX2 U1309 ( .A(n1176), .Z(n1238) );
  HS65_GS_FA1X4 U1310 ( .A0(n1179), .B0(n1178), .CI(n1177), .CO(n1174), .S0(
        n1180) );
  HS65_GS_IVX2 U1311 ( .A(n1180), .Z(n1234) );
  HS65_GS_FA1X4 U1312 ( .A0(n1183), .B0(n1182), .CI(n1181), .CO(n1178), .S0(
        n1184) );
  HS65_GS_IVX2 U1313 ( .A(n1184), .Z(n1230) );
  HS65_GS_FA1X4 U1314 ( .A0(n1187), .B0(n1186), .CI(n1185), .CO(n1182), .S0(
        n1188) );
  HS65_GS_IVX2 U1315 ( .A(n1188), .Z(n1226) );
  HS65_GS_FA1X4 U1316 ( .A0(n1191), .B0(n1190), .CI(n1189), .CO(n1186), .S0(
        n1192) );
  HS65_GS_IVX2 U1317 ( .A(n1192), .Z(n1222) );
  HS65_GS_FA1X4 U1318 ( .A0(n1195), .B0(n1194), .CI(n1193), .CO(n1190), .S0(
        n1196) );
  HS65_GS_IVX2 U1319 ( .A(n1196), .Z(n1218) );
  HS65_GS_FA1X4 U1320 ( .A0(n1199), .B0(n1198), .CI(n1197), .CO(n1194), .S0(
        n1200) );
  HS65_GS_IVX2 U1321 ( .A(n1200), .Z(n1214) );
  HS65_GS_FA1X4 U1322 ( .A0(n1203), .B0(n1202), .CI(n1201), .CO(n1198), .S0(
        n1204) );
  HS65_GS_IVX2 U1323 ( .A(n1204), .Z(n1209) );
  HS65_GS_FA1X4 U1324 ( .A0(p_b2[1]), .B0(n1206), .CI(n1205), .CO(n1202), .S0(
        n1207) );
  HS65_GS_IVX2 U1325 ( .A(n1207), .Z(n1211) );
  HS65_GS_FA1X4 U1326 ( .A0(p_b2[0]), .B0(p_b0[0]), .CI(p_b1[0]), .CO(n1205), 
        .S0(n1208) );
  HS65_GS_IVX2 U1327 ( .A(n1208), .Z(n1383) );
  HS65_GS_NAND2X2 U1328 ( .A(n1286), .B(p_a1[1]), .Z(n1285) );
  HS65_GS_NAND3AX3 U1329 ( .A(n1285), .B(p_a2[1]), .C(n1211), .Z(n1213) );
  HS65_GS_FA1X4 U1330 ( .A0(p_a2[2]), .B0(p_a1[2]), .CI(n1209), .CO(n1216), 
        .S0(n1290) );
  HS65_GS_FA1X4 U1331 ( .A0(p_a2[1]), .B0(n1211), .CI(n1210), .CO(n1212), .S0(
        n1286) );
  HS65_GS_CB4I1X4 U1332 ( .A(p_a1[1]), .B(n1286), .C(n1212), .D(n1213), .Z(
        n1289) );
  HS65_GS_NAND2X2 U1333 ( .A(n1290), .B(n1289), .Z(n1288) );
  HS65_GS_NAND2X2 U1334 ( .A(n1213), .B(n1288), .Z(n1215) );
  HS65_GS_NAND2X2 U1335 ( .A(n1216), .B(n1215), .Z(n1217) );
  HS65_GS_FA1X4 U1336 ( .A0(p_a2[3]), .B0(p_a1[3]), .CI(n1214), .CO(n1219), 
        .S0(n1294) );
  HS65_GSS_XOR2X3 U1337 ( .A(n1216), .B(n1215), .Z(n1293) );
  HS65_GS_NAND2X2 U1338 ( .A(n1294), .B(n1293), .Z(n1292) );
  HS65_GS_NAND2X2 U1339 ( .A(n1217), .B(n1292), .Z(n1220) );
  HS65_GS_NAND2X2 U1340 ( .A(n1219), .B(n1220), .Z(n1221) );
  HS65_GS_FA1X4 U1341 ( .A0(p_a2[4]), .B0(p_a1[4]), .CI(n1218), .CO(n1223), 
        .S0(n1298) );
  HS65_GSS_XOR2X3 U1342 ( .A(n1220), .B(n1219), .Z(n1297) );
  HS65_GS_NAND2X2 U1343 ( .A(n1298), .B(n1297), .Z(n1296) );
  HS65_GS_NAND2X2 U1344 ( .A(n1221), .B(n1296), .Z(n1224) );
  HS65_GS_NAND2X2 U1345 ( .A(n1223), .B(n1224), .Z(n1225) );
  HS65_GS_FA1X4 U1346 ( .A0(p_a2[5]), .B0(p_a1[5]), .CI(n1222), .CO(n1227), 
        .S0(n1302) );
  HS65_GSS_XOR2X3 U1347 ( .A(n1224), .B(n1223), .Z(n1301) );
  HS65_GS_NAND2X2 U1348 ( .A(n1302), .B(n1301), .Z(n1300) );
  HS65_GS_NAND2X2 U1349 ( .A(n1225), .B(n1300), .Z(n1228) );
  HS65_GS_NAND2X2 U1350 ( .A(n1227), .B(n1228), .Z(n1229) );
  HS65_GS_FA1X4 U1351 ( .A0(p_a2[6]), .B0(p_a1[6]), .CI(n1226), .CO(n1231), 
        .S0(n1306) );
  HS65_GSS_XOR2X3 U1352 ( .A(n1228), .B(n1227), .Z(n1305) );
  HS65_GS_NAND2X2 U1353 ( .A(n1306), .B(n1305), .Z(n1304) );
  HS65_GS_NAND2X2 U1354 ( .A(n1229), .B(n1304), .Z(n1232) );
  HS65_GS_NAND2X2 U1355 ( .A(n1231), .B(n1232), .Z(n1233) );
  HS65_GS_FA1X4 U1356 ( .A0(p_a2[7]), .B0(p_a1[7]), .CI(n1230), .CO(n1235), 
        .S0(n1310) );
  HS65_GSS_XOR2X3 U1357 ( .A(n1232), .B(n1231), .Z(n1309) );
  HS65_GS_NAND2X2 U1358 ( .A(n1310), .B(n1309), .Z(n1308) );
  HS65_GS_NAND2X2 U1359 ( .A(n1233), .B(n1308), .Z(n1236) );
  HS65_GS_NAND2X2 U1360 ( .A(n1235), .B(n1236), .Z(n1237) );
  HS65_GS_FA1X4 U1361 ( .A0(p_a2[8]), .B0(p_a1[8]), .CI(n1234), .CO(n1239), 
        .S0(n1314) );
  HS65_GSS_XOR2X3 U1362 ( .A(n1236), .B(n1235), .Z(n1313) );
  HS65_GS_NAND2X2 U1363 ( .A(n1314), .B(n1313), .Z(n1312) );
  HS65_GS_NAND2X2 U1364 ( .A(n1237), .B(n1312), .Z(n1240) );
  HS65_GS_NAND2X2 U1365 ( .A(n1239), .B(n1240), .Z(n1241) );
  HS65_GS_FA1X4 U1366 ( .A0(p_a2[9]), .B0(p_a1[9]), .CI(n1238), .CO(n1243), 
        .S0(n1318) );
  HS65_GSS_XOR2X3 U1367 ( .A(n1240), .B(n1239), .Z(n1317) );
  HS65_GS_NAND2X2 U1368 ( .A(n1318), .B(n1317), .Z(n1316) );
  HS65_GS_NAND2X2 U1369 ( .A(n1241), .B(n1316), .Z(n1244) );
  HS65_GS_NAND2X2 U1370 ( .A(n1243), .B(n1244), .Z(n1245) );
  HS65_GS_FA1X4 U1371 ( .A0(p_a2[10]), .B0(p_a1[10]), .CI(n1242), .CO(n1247), 
        .S0(n1322) );
  HS65_GSS_XOR2X3 U1372 ( .A(n1244), .B(n1243), .Z(n1321) );
  HS65_GS_NAND2X2 U1373 ( .A(n1322), .B(n1321), .Z(n1320) );
  HS65_GS_NAND2X2 U1374 ( .A(n1245), .B(n1320), .Z(n1248) );
  HS65_GS_NAND2X2 U1375 ( .A(n1247), .B(n1248), .Z(n1249) );
  HS65_GS_FA1X4 U1376 ( .A0(p_a2[11]), .B0(p_a1[11]), .CI(n1246), .CO(n1328), 
        .S0(n1326) );
  HS65_GSS_XOR2X3 U1377 ( .A(n1248), .B(n1247), .Z(n1325) );
  HS65_GS_NAND2X2 U1378 ( .A(n1326), .B(n1325), .Z(n1324) );
  HS65_GS_NAND2X2 U1379 ( .A(n1249), .B(n1324), .Z(n1329) );
  HS65_GS_PAO2X4 U1380 ( .A(n1328), .B(n1331), .P(n1329), .Z(n1251) );
  HS65_GS_FA1X4 U1381 ( .A0(p_a2[12]), .B0(p_a1[12]), .CI(n1250), .CO(n1252), 
        .S0(n1331) );
  HS65_GSS_XOR2X3 U1382 ( .A(n1251), .B(n1252), .Z(n1338) );
  HS65_GS_AO22X4 U1383 ( .A(n1337), .B(n1338), .C(n1252), .D(n1251), .Z(n1343)
         );
  HS65_GS_FA1X4 U1384 ( .A0(p_a1[13]), .B0(p_a2[13]), .CI(n1253), .CO(n1342), 
        .S0(n1337) );
  HS65_GS_FA1X4 U1385 ( .A0(p_b0[13]), .B0(p_b1[13]), .CI(p_b2[13]), .CO(n1261), .S0(n1254) );
  HS65_GS_FA1X4 U1386 ( .A0(n1256), .B0(n1255), .CI(n1254), .CO(n1260), .S0(
        n1160) );
  HS65_GS_IVX2 U1387 ( .A(n1257), .Z(n1258) );
  HS65_GS_FA1X4 U1388 ( .A0(p_a1[14]), .B0(p_a2[14]), .CI(n1258), .CO(n1267), 
        .S0(n1341) );
  HS65_GS_FA1X4 U1389 ( .A0(p_b0[14]), .B0(p_b1[14]), .CI(p_b2[14]), .CO(n1271), .S0(n1259) );
  HS65_GS_FA1X4 U1390 ( .A0(n1261), .B0(n1260), .CI(n1259), .CO(n1270), .S0(
        n1257) );
  HS65_GS_IVX2 U1391 ( .A(p_b0[15]), .Z(n1272) );
  HS65_GS_NAND2X2 U1392 ( .A(p_b2[15]), .B(p_b1[15]), .Z(n1273) );
  HS65_GS_OAI21X2 U1393 ( .A(p_b2[15]), .B(p_b1[15]), .C(n1273), .Z(n1262) );
  HS65_GS_MUXI21X2 U1394 ( .D0(p_b0[15]), .D1(n1272), .S0(n1262), .Z(n1269) );
  HS65_GS_IVX2 U1395 ( .A(n1263), .Z(n1266) );
  HS65_GS_IVX2 U1396 ( .A(n1264), .Z(n1283) );
  HS65_GS_FA1X4 U1397 ( .A0(p_a1[15]), .B0(p_a2[15]), .CI(n1265), .CO(n1277), 
        .S0(n1263) );
  HS65_GS_FA1X4 U1398 ( .A0(n1268), .B0(n1267), .CI(n1266), .CO(n1279), .S0(
        n1264) );
  HS65_GS_FA1X4 U1399 ( .A0(n1271), .B0(n1270), .CI(n1269), .CO(n1275), .S0(
        n1265) );
  HS65_GS_OAI32X2 U1400 ( .A(p_b0[15]), .B(p_b2[15]), .C(p_b1[15]), .D(n1273), 
        .E(n1272), .Z(n1274) );
  HS65_GSS_XNOR2X3 U1401 ( .A(n1275), .B(n1274), .Z(n1278) );
  HS65_GSS_XNOR2X3 U1402 ( .A(n1279), .B(n1278), .Z(n1276) );
  HS65_GS_NOR2X2 U1403 ( .A(n1277), .B(n1276), .Z(n1280) );
  HS65_GS_AND2X4 U1404 ( .A(n1277), .B(n1276), .Z(n1284) );
  HS65_GS_OA12X4 U1405 ( .A(n1280), .B(n1284), .C(valid_T3), .Z(n1282) );
  HS65_GS_NAND2X2 U1406 ( .A(n1279), .B(n1278), .Z(n1281) );
  HS65_GS_NOR3AX2 U1407 ( .A(n1281), .B(n1784), .C(n1280), .Z(n1782) );
  HS65_GS_AOI12X2 U1408 ( .A(n1283), .B(n1282), .C(n1782), .Z(n1387) );
  HS65_GS_IVX2 U1409 ( .A(n1387), .Z(n1335) );
  HS65_GS_OAI12X3 U1410 ( .A(n1284), .B(n1283), .C(n1782), .Z(n1344) );
  HS65_GS_OAI112X1 U1411 ( .A(n1286), .B(p_a1[1]), .C(n1344), .D(n1285), .Z(
        n1287) );
  HS65_GS_AO22X4 U1412 ( .A(data_out[1]), .B(n1784), .C(n1335), .D(n1287), .Z(
        n1883) );
  HS65_GS_MUXI21X2 U1413 ( .D0(n1534), .D1(n1661), .S0(valid_in), .Z(n1882) );
  HS65_GS_OAI112X1 U1414 ( .A(n1290), .B(n1289), .C(n1344), .D(n1288), .Z(
        n1291) );
  HS65_GS_AO22X4 U1415 ( .A(data_out[2]), .B(n1784), .C(n1335), .D(n1291), .Z(
        n1880) );
  HS65_GS_MUXI21X2 U1416 ( .D0(n1532), .D1(n1659), .S0(n1366), .Z(n1879) );
  HS65_GS_OAI112X1 U1417 ( .A(n1294), .B(n1293), .C(n1344), .D(n1292), .Z(
        n1295) );
  HS65_GS_AO22X4 U1418 ( .A(data_out[3]), .B(n1784), .C(n1335), .D(n1295), .Z(
        n1877) );
  HS65_GS_MUXI21X2 U1419 ( .D0(n1530), .D1(n1657), .S0(n1792), .Z(n1876) );
  HS65_GS_OAI112X1 U1420 ( .A(n1298), .B(n1297), .C(n1344), .D(n1296), .Z(
        n1299) );
  HS65_GS_AO22X4 U1421 ( .A(data_out[4]), .B(n1784), .C(n1335), .D(n1299), .Z(
        n1874) );
  HS65_GS_BFX4 U1422 ( .A(n1366), .Z(n1361) );
  HS65_GS_MUXI21X2 U1423 ( .D0(n1528), .D1(n1655), .S0(n1361), .Z(n1873) );
  HS65_GS_OAI112X1 U1424 ( .A(n1302), .B(n1301), .C(n1344), .D(n1300), .Z(
        n1303) );
  HS65_GS_AO22X4 U1425 ( .A(data_out[5]), .B(n1784), .C(n1335), .D(n1303), .Z(
        n1871) );
  HS65_GS_MUXI21X2 U1426 ( .D0(n1526), .D1(n1653), .S0(n1361), .Z(n1870) );
  HS65_GS_OAI112X1 U1427 ( .A(n1306), .B(n1305), .C(n1344), .D(n1304), .Z(
        n1307) );
  HS65_GS_AO22X4 U1428 ( .A(data_out[6]), .B(n1784), .C(n1335), .D(n1307), .Z(
        n1868) );
  HS65_GS_MUXI21X2 U1429 ( .D0(n1524), .D1(n1651), .S0(n1361), .Z(n1867) );
  HS65_GS_OAI112X1 U1430 ( .A(n1310), .B(n1309), .C(n1344), .D(n1308), .Z(
        n1311) );
  HS65_GS_AO22X4 U1431 ( .A(data_out[7]), .B(n1784), .C(n1335), .D(n1311), .Z(
        n1865) );
  HS65_GS_MUXI21X2 U1432 ( .D0(n1522), .D1(n1649), .S0(n1361), .Z(n1864) );
  HS65_GS_OAI112X1 U1433 ( .A(n1314), .B(n1313), .C(n1344), .D(n1312), .Z(
        n1315) );
  HS65_GS_AO22X4 U1434 ( .A(data_out[8]), .B(n1784), .C(n1335), .D(n1315), .Z(
        n1862) );
  HS65_GS_MUXI21X2 U1435 ( .D0(n1520), .D1(n1647), .S0(n1361), .Z(n1861) );
  HS65_GS_OAI112X1 U1436 ( .A(n1318), .B(n1317), .C(n1344), .D(n1316), .Z(
        n1319) );
  HS65_GS_AO22X4 U1437 ( .A(data_out[9]), .B(n1784), .C(n1335), .D(n1319), .Z(
        n1859) );
  HS65_GS_MUXI21X2 U1438 ( .D0(n1518), .D1(n1645), .S0(n1361), .Z(n1858) );
  HS65_GS_OAI112X1 U1439 ( .A(n1322), .B(n1321), .C(n1344), .D(n1320), .Z(
        n1323) );
  HS65_GS_AO22X4 U1440 ( .A(data_out[10]), .B(n1784), .C(n1335), .D(n1323), 
        .Z(n1856) );
  HS65_GS_MUXI21X2 U1441 ( .D0(n1516), .D1(n1643), .S0(n1382), .Z(n1855) );
  HS65_GS_OAI112X1 U1442 ( .A(n1326), .B(n1325), .C(n1344), .D(n1324), .Z(
        n1327) );
  HS65_GS_AO22X4 U1443 ( .A(data_out[11]), .B(n1784), .C(n1335), .D(n1327), 
        .Z(n1853) );
  HS65_GS_MUXI21X2 U1444 ( .D0(n1514), .D1(n1641), .S0(n1361), .Z(n1852) );
  HS65_GS_IVX2 U1445 ( .A(data_out[12]), .Z(n1334) );
  HS65_GS_MUXI21X2 U1446 ( .D0(n1641), .D1(n1334), .S0(n1382), .Z(n1851) );
  HS65_GSS_XOR2X3 U1447 ( .A(n1329), .B(n1328), .Z(n1332) );
  HS65_GS_OAI21X2 U1448 ( .A(n1331), .B(n1332), .C(n1344), .Z(n1330) );
  HS65_GS_CBI4I1X3 U1449 ( .A(n1332), .B(n1331), .C(n1330), .D(n1335), .Z(
        n1333) );
  HS65_GS_OAI21X2 U1450 ( .A(valid_T3), .B(n1334), .C(n1333), .Z(n1850) );
  HS65_GS_MUXI21X2 U1451 ( .D0(n1512), .D1(n1639), .S0(n1382), .Z(n1849) );
  HS65_GS_IVX2 U1452 ( .A(data_out[13]), .Z(n1340) );
  HS65_GS_MUXI21X2 U1453 ( .D0(n1639), .D1(n1340), .S0(n1382), .Z(n1848) );
  HS65_GS_OAI21X2 U1454 ( .A(n1337), .B(n1338), .C(n1344), .Z(n1336) );
  HS65_GS_CBI4I1X3 U1455 ( .A(n1338), .B(n1337), .C(n1336), .D(n1335), .Z(
        n1339) );
  HS65_GS_OAI21X2 U1456 ( .A(valid_T3), .B(n1340), .C(n1339), .Z(n1847) );
  HS65_GS_MUXI21X2 U1457 ( .D0(n1510), .D1(n1637), .S0(n1382), .Z(n1846) );
  HS65_GS_FA1X4 U1458 ( .A0(n1343), .B0(n1342), .CI(n1341), .CO(n1268), .S0(
        n1346) );
  HS65_GS_IVX2 U1459 ( .A(n1344), .Z(n1384) );
  HS65_GS_AOI12X2 U1460 ( .A(data_out[14]), .B(n1784), .C(n1384), .Z(n1345) );
  HS65_GS_OAI21X2 U1461 ( .A(n1387), .B(n1346), .C(n1345), .Z(n1844) );
  HS65_GS_MUXI21X2 U1462 ( .D0(n1710), .D1(n1635), .S0(n1382), .Z(n1843) );
  HS65_GS_IVX2 U1463 ( .A(data_out[15]), .Z(n1783) );
  HS65_GS_MUXI21X2 U1464 ( .D0(n1635), .D1(n1783), .S0(n1382), .Z(n1842) );
  HS65_GS_MUXI21X2 U1465 ( .D0(n1677), .D1(n1347), .S0(valid_in), .Z(n1840) );
  HS65_GS_MUXI21X2 U1466 ( .D0(n1347), .D1(n1348), .S0(valid_in), .Z(n1839) );
  HS65_GS_MUXI21X2 U1467 ( .D0(n1714), .D1(n1349), .S0(n1366), .Z(n1838) );
  HS65_GS_MUXI21X2 U1468 ( .D0(n1349), .D1(n1350), .S0(valid_in), .Z(n1837) );
  HS65_GS_MUX21X4 U1469 ( .D0(x_reg2[2]), .D1(x_z2[2]), .S0(n1792), .Z(n1836)
         );
  HS65_GS_MUXI21X2 U1470 ( .D0(n1706), .D1(n1351), .S0(valid_in), .Z(n1835) );
  HS65_GS_MUX21X4 U1471 ( .D0(x_reg2[3]), .D1(x_z2[3]), .S0(n1366), .Z(n1834)
         );
  HS65_GS_MUXI21X2 U1472 ( .D0(n1704), .D1(n1352), .S0(n1792), .Z(n1833) );
  HS65_GS_MUX21X4 U1473 ( .D0(x_reg2[4]), .D1(x_z2[4]), .S0(n1366), .Z(n1832)
         );
  HS65_GS_MUXI21X2 U1474 ( .D0(n1702), .D1(n1353), .S0(valid_in), .Z(n1831) );
  HS65_GS_MUX21X4 U1475 ( .D0(x_reg2[5]), .D1(x_z2[5]), .S0(n1366), .Z(n1830)
         );
  HS65_GS_MUXI21X2 U1476 ( .D0(n1700), .D1(n1354), .S0(n1366), .Z(n1829) );
  HS65_GS_MUX21X4 U1477 ( .D0(x_reg2[6]), .D1(x_z2[6]), .S0(n1366), .Z(n1828)
         );
  HS65_GS_MUXI21X2 U1478 ( .D0(n1698), .D1(n1355), .S0(n1361), .Z(n1827) );
  HS65_GS_MUX21X4 U1479 ( .D0(x_reg2[7]), .D1(x_z2[7]), .S0(n1792), .Z(n1826)
         );
  HS65_GS_MUXI21X2 U1480 ( .D0(n1696), .D1(n1356), .S0(n1361), .Z(n1825) );
  HS65_GS_MUX21X4 U1481 ( .D0(x_reg2[8]), .D1(x_z2[8]), .S0(valid_in), .Z(
        n1824) );
  HS65_GS_MUXI21X2 U1482 ( .D0(n1694), .D1(n1357), .S0(n1361), .Z(n1823) );
  HS65_GS_MUX21X4 U1483 ( .D0(x_reg2[9]), .D1(x_z2[9]), .S0(n1366), .Z(n1822)
         );
  HS65_GS_MUXI21X2 U1484 ( .D0(n1692), .D1(n1358), .S0(n1361), .Z(n1821) );
  HS65_GS_MUX21X4 U1485 ( .D0(x_reg2[10]), .D1(x_z2[10]), .S0(n1792), .Z(n1820) );
  HS65_GS_MUXI21X2 U1486 ( .D0(n1690), .D1(n1359), .S0(n1361), .Z(n1819) );
  HS65_GS_MUX21X4 U1487 ( .D0(x_reg2[11]), .D1(x_z2[11]), .S0(n1792), .Z(n1818) );
  HS65_GS_MUXI21X2 U1488 ( .D0(n1688), .D1(n1360), .S0(n1382), .Z(n1817) );
  HS65_GS_MUX21X4 U1489 ( .D0(x_reg2[12]), .D1(x_z2[12]), .S0(valid_in), .Z(
        n1816) );
  HS65_GS_MUXI21X2 U1490 ( .D0(n1686), .D1(n1362), .S0(n1361), .Z(n1815) );
  HS65_GS_MUX21X4 U1491 ( .D0(x_reg2[13]), .D1(x_z2[13]), .S0(n1366), .Z(n1814) );
  HS65_GS_MUXI21X2 U1492 ( .D0(n1684), .D1(n1363), .S0(n1382), .Z(n1813) );
  HS65_GS_MUX21X4 U1493 ( .D0(x_reg2[14]), .D1(x_z2[14]), .S0(valid_in), .Z(
        n1812) );
  HS65_GS_MUXI21X2 U1494 ( .D0(n1682), .D1(n1364), .S0(n1382), .Z(n1811) );
  HS65_GS_MUXI21X2 U1495 ( .D0(n1727), .D1(n1680), .S0(n1382), .Z(n1810) );
  HS65_GS_MUXI21X2 U1496 ( .D0(n1680), .D1(n1365), .S0(n1382), .Z(n1809) );
  HS65_GS_MUX21X4 U1497 ( .D0(x_z1[0]), .D1(data_in[0]), .S0(n1792), .Z(n1808)
         );
  HS65_GS_MUX21X4 U1498 ( .D0(x_z1[1]), .D1(data_in[1]), .S0(n1366), .Z(n1807)
         );
  HS65_GS_MUX21X4 U1499 ( .D0(x_z1[2]), .D1(data_in[2]), .S0(n1792), .Z(n1806)
         );
  HS65_GS_MUX21X4 U1500 ( .D0(x_z1[3]), .D1(data_in[3]), .S0(n1366), .Z(n1805)
         );
  HS65_GS_MUX21X4 U1501 ( .D0(x_z1[4]), .D1(data_in[4]), .S0(n1366), .Z(n1804)
         );
  HS65_GS_MUX21X4 U1502 ( .D0(x_z1[5]), .D1(data_in[5]), .S0(valid_in), .Z(
        n1803) );
  HS65_GS_MUX21X4 U1503 ( .D0(x_z1[6]), .D1(data_in[6]), .S0(valid_in), .Z(
        n1802) );
  HS65_GS_MUX21X4 U1504 ( .D0(x_z1[7]), .D1(data_in[7]), .S0(valid_in), .Z(
        n1801) );
  HS65_GS_MUX21X4 U1505 ( .D0(x_z1[8]), .D1(data_in[8]), .S0(n1366), .Z(n1800)
         );
  HS65_GS_MUX21X4 U1506 ( .D0(x_z1[9]), .D1(data_in[9]), .S0(n1792), .Z(n1799)
         );
  HS65_GS_MUX21X4 U1507 ( .D0(x_z1[10]), .D1(data_in[10]), .S0(valid_in), .Z(
        n1798) );
  HS65_GS_MUX21X4 U1508 ( .D0(x_z1[11]), .D1(data_in[11]), .S0(n1366), .Z(
        n1797) );
  HS65_GS_MUX21X4 U1509 ( .D0(x_z1[12]), .D1(data_in[12]), .S0(valid_in), .Z(
        n1796) );
  HS65_GS_MUX21X4 U1510 ( .D0(x_z1[13]), .D1(data_in[13]), .S0(valid_in), .Z(
        n1795) );
  HS65_GS_MUX21X4 U1511 ( .D0(x_z1[14]), .D1(data_in[14]), .S0(n1792), .Z(
        n1794) );
  HS65_GSS_XNOR2X3 U1512 ( .A(y_z2[15]), .B(n1367), .Z(n1511) );
  HS65_GS_AND2X4 U1513 ( .A(n1511), .B(y_z2[14]), .Z(\mul_a2/fa1_c2[28] ) );
  HS65_GS_HA1X4 U1514 ( .A0(n1710), .B0(n1368), .CO(n1367), .S0(n1513) );
  HS65_GS_AND2X4 U1515 ( .A(n1513), .B(y_z2[13]), .Z(\mul_a2/fa1_c2[27] ) );
  HS65_GS_HA1X4 U1516 ( .A0(n1510), .B0(n1369), .CO(n1368), .S0(n1515) );
  HS65_GS_AND2X4 U1517 ( .A(n1515), .B(y_z2[12]), .Z(\mul_a2/fa1_c2[26] ) );
  HS65_GS_HA1X4 U1518 ( .A0(n1512), .B0(n1370), .CO(n1369), .S0(n1517) );
  HS65_GS_AND2X4 U1519 ( .A(n1517), .B(y_z2[11]), .Z(\mul_a2/fa1_c2[25] ) );
  HS65_GS_HA1X4 U1520 ( .A0(n1514), .B0(n1371), .CO(n1370), .S0(n1519) );
  HS65_GS_AND2X4 U1521 ( .A(y_z2[10]), .B(n1519), .Z(\mul_a2/fa1_c2[24] ) );
  HS65_GS_HA1X4 U1522 ( .A0(n1516), .B0(n1372), .CO(n1371), .S0(n1521) );
  HS65_GS_AND2X4 U1523 ( .A(y_z2[9]), .B(n1521), .Z(\mul_a2/fa1_c2[23] ) );
  HS65_GS_HA1X4 U1524 ( .A0(n1518), .B0(n1373), .CO(n1372), .S0(n1523) );
  HS65_GS_AND2X4 U1525 ( .A(n1523), .B(y_z2[8]), .Z(\mul_a2/fa1_c2[22] ) );
  HS65_GS_HA1X4 U1526 ( .A0(n1520), .B0(n1374), .CO(n1373), .S0(n1525) );
  HS65_GS_AND2X4 U1527 ( .A(y_z2[7]), .B(n1525), .Z(\mul_a2/fa1_c2[21] ) );
  HS65_GS_HA1X4 U1528 ( .A0(n1522), .B0(n1375), .CO(n1374), .S0(n1527) );
  HS65_GS_AND2X4 U1529 ( .A(y_z2[6]), .B(n1527), .Z(\mul_a2/fa1_c2[20] ) );
  HS65_GS_HA1X4 U1530 ( .A0(n1524), .B0(n1376), .CO(n1375), .S0(n1529) );
  HS65_GS_AND2X4 U1531 ( .A(y_z2[5]), .B(n1529), .Z(\mul_a2/fa1_c2[19] ) );
  HS65_GS_HA1X4 U1532 ( .A0(n1526), .B0(n1377), .CO(n1376), .S0(n1531) );
  HS65_GS_AND2X4 U1533 ( .A(n1531), .B(y_z2[4]), .Z(\mul_a2/fa1_c2[18] ) );
  HS65_GS_HA1X4 U1534 ( .A0(n1528), .B0(n1378), .CO(n1377), .S0(n1533) );
  HS65_GS_AND2X4 U1535 ( .A(n1533), .B(y_z2[3]), .Z(\mul_a2/fa1_c2[17] ) );
  HS65_GS_HA1X4 U1536 ( .A0(n1530), .B0(n1379), .CO(n1378), .S0(n1535) );
  HS65_GS_AND2X4 U1537 ( .A(n1535), .B(y_z2[2]), .Z(\mul_a2/fa1_c2[16] ) );
  HS65_GS_HA1X4 U1538 ( .A0(n1532), .B0(n1380), .CO(n1379), .S0(n1536) );
  HS65_GS_AND2X4 U1539 ( .A(n1536), .B(y_z2[1]), .Z(\mul_a2/fa1_c2[15] ) );
  HS65_GS_HA1X4 U1540 ( .A0(n1534), .B0(n1381), .CO(n1380), .S0(n1537) );
  HS65_GS_AND2X4 U1541 ( .A(y_z2[0]), .B(n1537), .Z(\mul_a2/fa1_c2[14] ) );
  HS65_GS_MUXI21X2 U1542 ( .D0(n1707), .D1(n1712), .S0(n1382), .Z(n1888) );
  HS65_GS_FA1X4 U1543 ( .A0(p_a2[0]), .B0(p_a1[0]), .CI(n1383), .CO(n1210), 
        .S0(n1386) );
  HS65_GS_AOI12X2 U1544 ( .A(data_out[0]), .B(n1784), .C(n1384), .Z(n1385) );
  HS65_GS_OAI21X2 U1545 ( .A(n1387), .B(n1386), .C(n1385), .Z(n1886) );
  HS65_GS_MUXI21X2 U1546 ( .D0(n1708), .D1(n1713), .S0(n1792), .Z(n1885) );
  HS65_GS_HA1X4 U1547 ( .A0(n1637), .B0(n1388), .CO(n1431), .S0(n1620) );
  HS65_GS_AND2X4 U1548 ( .A(n1620), .B(y_z1[12]), .Z(\mul_a1/fa1_c0[15] ) );
  HS65_GS_HA1X4 U1549 ( .A0(n1639), .B0(n1389), .CO(n1388), .S0(n1621) );
  HS65_GS_AND2X4 U1550 ( .A(n1621), .B(y_z1[11]), .Z(\mul_a1/fa1_c0[14] ) );
  HS65_GS_HA1X4 U1551 ( .A0(n1641), .B0(n1390), .CO(n1389), .S0(n1622) );
  HS65_GS_AND2X4 U1552 ( .A(n1622), .B(y_z1[10]), .Z(\mul_a1/fa1_c0[13] ) );
  HS65_GS_HA1X4 U1553 ( .A0(n1643), .B0(n1391), .CO(n1390), .S0(n1623) );
  HS65_GS_AND2X4 U1554 ( .A(n1623), .B(y_z1[9]), .Z(\mul_a1/fa1_c0[12] ) );
  HS65_GS_HA1X4 U1555 ( .A0(n1645), .B0(n1392), .CO(n1391), .S0(n1624) );
  HS65_GS_AND2X4 U1556 ( .A(n1624), .B(y_z1[8]), .Z(\mul_a1/fa1_c0[11] ) );
  HS65_GS_HA1X4 U1557 ( .A0(n1647), .B0(n1393), .CO(n1392), .S0(n1625) );
  HS65_GS_AND2X4 U1558 ( .A(n1625), .B(y_z1[7]), .Z(\mul_a1/fa1_c0[10] ) );
  HS65_GS_HA1X4 U1559 ( .A0(n1649), .B0(n1394), .CO(n1393), .S0(n1626) );
  HS65_GS_AND2X4 U1560 ( .A(n1626), .B(y_z1[6]), .Z(\mul_a1/fa1_c0[9] ) );
  HS65_GS_HA1X4 U1561 ( .A0(n1651), .B0(n1395), .CO(n1394), .S0(n1627) );
  HS65_GS_AND2X4 U1562 ( .A(n1627), .B(y_z1[5]), .Z(\mul_a1/fa1_c0[8] ) );
  HS65_GS_HA1X4 U1563 ( .A0(n1653), .B0(n1396), .CO(n1395), .S0(n1628) );
  HS65_GS_AND2X4 U1564 ( .A(n1628), .B(y_z1[4]), .Z(\mul_a1/fa1_c0[7] ) );
  HS65_GS_HA1X4 U1565 ( .A0(n1655), .B0(n1397), .CO(n1396), .S0(n1629) );
  HS65_GS_AND2X4 U1566 ( .A(n1629), .B(y_z1[3]), .Z(\mul_a1/fa1_c0[6] ) );
  HS65_GS_HA1X4 U1567 ( .A0(n1657), .B0(n1398), .CO(n1397), .S0(n1630) );
  HS65_GS_AND2X4 U1568 ( .A(n1630), .B(y_z1[2]), .Z(\mul_a1/fa1_c0[5] ) );
  HS65_GS_HA1X4 U1569 ( .A0(n1659), .B0(n1399), .CO(n1398), .S0(n1631) );
  HS65_GS_AND2X4 U1570 ( .A(n1631), .B(y_z1[1]), .Z(\mul_a1/fa1_c0[4] ) );
  HS65_GS_HA1X4 U1571 ( .A0(n1661), .B0(n1400), .CO(n1399), .S0(n1401) );
  HS65_GS_AND2X4 U1572 ( .A(n1401), .B(y_z1[0]), .Z(\mul_a1/fa1_c0[3] ) );
  HS65_GSS_XNOR2X3 U1573 ( .A(y_z1[15]), .B(n1402), .Z(n1417) );
  HS65_GSS_XNOR2X3 U1574 ( .A(n1417), .B(n1639), .Z(\mul_a1/fa1_s1[24] ) );
  HS65_GS_HA1X4 U1575 ( .A0(n1637), .B0(n1403), .CO(n1402), .S0(n1418) );
  HS65_GSS_XNOR2X3 U1576 ( .A(n1418), .B(n1641), .Z(\mul_a1/fa1_s1[23] ) );
  HS65_GS_HA1X4 U1577 ( .A0(n1639), .B0(n1404), .CO(n1403), .S0(n1419) );
  HS65_GSS_XNOR2X3 U1578 ( .A(n1419), .B(n1643), .Z(\mul_a1/fa1_s1[22] ) );
  HS65_GS_HA1X4 U1579 ( .A0(n1641), .B0(n1405), .CO(n1404), .S0(n1420) );
  HS65_GSS_XNOR2X3 U1580 ( .A(n1420), .B(n1645), .Z(\mul_a1/fa1_s1[21] ) );
  HS65_GS_HA1X4 U1581 ( .A0(n1643), .B0(n1406), .CO(n1405), .S0(n1421) );
  HS65_GSS_XNOR2X3 U1582 ( .A(n1421), .B(n1647), .Z(\mul_a1/fa1_s1[20] ) );
  HS65_GS_HA1X4 U1583 ( .A0(n1645), .B0(n1407), .CO(n1406), .S0(n1422) );
  HS65_GSS_XNOR2X3 U1584 ( .A(n1422), .B(n1649), .Z(\mul_a1/fa1_s1[19] ) );
  HS65_GS_HA1X4 U1585 ( .A0(n1647), .B0(n1408), .CO(n1407), .S0(n1423) );
  HS65_GSS_XNOR2X3 U1586 ( .A(n1423), .B(n1651), .Z(\mul_a1/fa1_s1[18] ) );
  HS65_GS_HA1X4 U1587 ( .A0(n1649), .B0(n1409), .CO(n1408), .S0(n1424) );
  HS65_GSS_XNOR2X3 U1588 ( .A(n1424), .B(n1653), .Z(\mul_a1/fa1_s1[17] ) );
  HS65_GS_HA1X4 U1589 ( .A0(n1651), .B0(n1410), .CO(n1409), .S0(n1425) );
  HS65_GSS_XNOR2X3 U1590 ( .A(n1425), .B(n1655), .Z(\mul_a1/fa1_s1[16] ) );
  HS65_GS_HA1X4 U1591 ( .A0(n1653), .B0(n1411), .CO(n1410), .S0(n1426) );
  HS65_GSS_XNOR2X3 U1592 ( .A(n1426), .B(n1657), .Z(\mul_a1/fa1_s1[15] ) );
  HS65_GS_HA1X4 U1593 ( .A0(n1655), .B0(n1412), .CO(n1411), .S0(n1427) );
  HS65_GSS_XNOR2X3 U1594 ( .A(n1427), .B(n1659), .Z(\mul_a1/fa1_s1[14] ) );
  HS65_GS_HA1X4 U1595 ( .A0(n1657), .B0(n1413), .CO(n1412), .S0(n1428) );
  HS65_GSS_XNOR2X3 U1596 ( .A(n1428), .B(n1661), .Z(\mul_a1/fa1_s1[13] ) );
  HS65_GS_HA1X4 U1597 ( .A0(n1659), .B0(n1414), .CO(n1413), .S0(n1429) );
  HS65_GSS_XNOR2X3 U1598 ( .A(n1429), .B(n1713), .Z(\mul_a1/fa1_s1[12] ) );
  HS65_GS_HA1X4 U1599 ( .A0(n1661), .B0(n1415), .CO(n1414), .S0(n1430) );
  HS65_GSS_XNOR2X3 U1600 ( .A(n1430), .B(n1712), .Z(\mul_a1/fa1_s1[11] ) );
  HS65_GS_AND2X4 U1601 ( .A(n1416), .B(y_z1[14]), .Z(\mul_a1/fa1_c1[25] ) );
  HS65_GS_AND2X4 U1602 ( .A(n1417), .B(y_z1[13]), .Z(\mul_a1/fa1_c1[24] ) );
  HS65_GS_AND2X4 U1603 ( .A(n1418), .B(y_z1[12]), .Z(\mul_a1/fa1_c1[23] ) );
  HS65_GS_AND2X4 U1604 ( .A(n1419), .B(y_z1[11]), .Z(\mul_a1/fa1_c1[22] ) );
  HS65_GS_AND2X4 U1605 ( .A(n1420), .B(y_z1[10]), .Z(\mul_a1/fa1_c1[21] ) );
  HS65_GS_AND2X4 U1606 ( .A(n1421), .B(y_z1[9]), .Z(\mul_a1/fa1_c1[20] ) );
  HS65_GS_AND2X4 U1607 ( .A(n1422), .B(y_z1[8]), .Z(\mul_a1/fa1_c1[19] ) );
  HS65_GS_AND2X4 U1608 ( .A(n1423), .B(y_z1[7]), .Z(\mul_a1/fa1_c1[18] ) );
  HS65_GS_AND2X4 U1609 ( .A(n1424), .B(y_z1[6]), .Z(\mul_a1/fa1_c1[17] ) );
  HS65_GS_AND2X4 U1610 ( .A(n1425), .B(y_z1[5]), .Z(\mul_a1/fa1_c1[16] ) );
  HS65_GS_AND2X4 U1611 ( .A(n1426), .B(y_z1[4]), .Z(\mul_a1/fa1_c1[15] ) );
  HS65_GS_AND2X4 U1612 ( .A(n1427), .B(y_z1[3]), .Z(\mul_a1/fa1_c1[14] ) );
  HS65_GS_AND2X4 U1613 ( .A(n1428), .B(y_z1[2]), .Z(\mul_a1/fa1_c1[13] ) );
  HS65_GS_AND2X4 U1614 ( .A(n1429), .B(y_z1[1]), .Z(\mul_a1/fa1_c1[12] ) );
  HS65_GS_AND2X4 U1615 ( .A(n1430), .B(y_z1[0]), .Z(\mul_a1/fa1_c1[11] ) );
  HS65_GSS_XNOR2X3 U1616 ( .A(y_z1[15]), .B(n1431), .Z(n1619) );
  HS65_GS_AND2X4 U1617 ( .A(n1619), .B(y_z1[13]), .Z(\mul_a1/fa1_c0[16] ) );
  HS65_GS_IVX2 U1618 ( .A(n1447), .Z(n1744) );
  HS65_GS_FA1X4 U1619 ( .A0(n1434), .B0(n1433), .CI(n1432), .CO(n951), .S0(
        n1435) );
  HS65_GS_OAI21X2 U1620 ( .A(n1744), .B(n1435), .C(n1745), .Z(
        \mul_a1/result_sat[14] ) );
  HS65_GS_FA1X4 U1621 ( .A0(n1438), .B0(n1437), .CI(n1436), .CO(n762), .S0(
        n1439) );
  HS65_GS_AO12X4 U1622 ( .A(n1439), .B(n1447), .C(n1449), .Z(
        \mul_a1/result_sat[11] ) );
  HS65_GS_FA1X4 U1623 ( .A0(n1442), .B0(n1441), .CI(n1440), .CO(n1436), .S0(
        n1443) );
  HS65_GS_OA12X4 U1624 ( .A(n1449), .B(n1443), .C(n1447), .Z(
        \mul_a1/result_sat[10] ) );
  HS65_GS_FA1X4 U1625 ( .A0(n1446), .B0(n1445), .CI(n1444), .CO(n1441), .S0(
        n1448) );
  HS65_GS_OA12X4 U1626 ( .A(n1449), .B(n1448), .C(n1447), .Z(
        \mul_a1/result_sat[9] ) );
  HS65_GS_OAI21X2 U1627 ( .A(n1452), .B(n1451), .C(n1450), .Z(n1453) );
  HS65_GS_OAI21X2 U1628 ( .A(n1744), .B(n1453), .C(n1745), .Z(
        \mul_a1/result_sat[1] ) );
  HS65_GS_HA1X4 U1629 ( .A0(n1510), .B0(n1454), .CO(n1709), .S0(n1482) );
  HS65_GSS_XNOR2X3 U1630 ( .A(y_z2[15]), .B(n1455), .Z(n1481) );
  HS65_GSS_XOR2X3 U1631 ( .A(n1482), .B(n1481), .Z(\mul_a2/fa1_s1[22] ) );
  HS65_GS_HA1X4 U1632 ( .A0(n1510), .B0(n1456), .CO(n1455), .S0(n1484) );
  HS65_GS_HA1X4 U1633 ( .A0(n1512), .B0(n1457), .CO(n1454), .S0(n1483) );
  HS65_GSS_XOR2X3 U1634 ( .A(n1484), .B(n1483), .Z(\mul_a2/fa1_s1[21] ) );
  HS65_GS_HA1X4 U1635 ( .A0(n1512), .B0(n1458), .CO(n1456), .S0(n1486) );
  HS65_GS_HA1X4 U1636 ( .A0(n1514), .B0(n1459), .CO(n1457), .S0(n1485) );
  HS65_GSS_XOR2X3 U1637 ( .A(n1486), .B(n1485), .Z(\mul_a2/fa1_s1[20] ) );
  HS65_GS_HA1X4 U1638 ( .A0(n1514), .B0(n1460), .CO(n1458), .S0(n1488) );
  HS65_GS_HA1X4 U1639 ( .A0(n1516), .B0(n1461), .CO(n1459), .S0(n1487) );
  HS65_GSS_XOR2X3 U1640 ( .A(n1488), .B(n1487), .Z(\mul_a2/fa1_s1[19] ) );
  HS65_GS_HA1X4 U1641 ( .A0(n1518), .B0(n1462), .CO(n1461), .S0(n1490) );
  HS65_GS_HA1X4 U1642 ( .A0(n1516), .B0(n1463), .CO(n1460), .S0(n1489) );
  HS65_GSS_XOR2X3 U1643 ( .A(n1490), .B(n1489), .Z(\mul_a2/fa1_s1[18] ) );
  HS65_GS_HA1X4 U1644 ( .A0(n1520), .B0(n1464), .CO(n1462), .S0(n1492) );
  HS65_GS_HA1X4 U1645 ( .A0(n1518), .B0(n1465), .CO(n1463), .S0(n1491) );
  HS65_GSS_XOR2X3 U1646 ( .A(n1492), .B(n1491), .Z(\mul_a2/fa1_s1[17] ) );
  HS65_GS_HA1X4 U1647 ( .A0(n1522), .B0(n1466), .CO(n1464), .S0(n1494) );
  HS65_GS_HA1X4 U1648 ( .A0(n1520), .B0(n1467), .CO(n1465), .S0(n1493) );
  HS65_GSS_XOR2X3 U1649 ( .A(n1494), .B(n1493), .Z(\mul_a2/fa1_s1[16] ) );
  HS65_GS_HA1X4 U1650 ( .A0(n1524), .B0(n1468), .CO(n1466), .S0(n1496) );
  HS65_GS_HA1X4 U1651 ( .A0(n1522), .B0(n1469), .CO(n1467), .S0(n1495) );
  HS65_GSS_XOR2X3 U1652 ( .A(n1496), .B(n1495), .Z(\mul_a2/fa1_s1[15] ) );
  HS65_GS_HA1X4 U1653 ( .A0(n1524), .B0(n1470), .CO(n1469), .S0(n1498) );
  HS65_GS_HA1X4 U1654 ( .A0(n1526), .B0(n1471), .CO(n1468), .S0(n1497) );
  HS65_GSS_XOR2X3 U1655 ( .A(n1498), .B(n1497), .Z(\mul_a2/fa1_s1[14] ) );
  HS65_GS_HA1X4 U1656 ( .A0(n1526), .B0(n1472), .CO(n1470), .S0(n1500) );
  HS65_GS_HA1X4 U1657 ( .A0(n1528), .B0(n1473), .CO(n1471), .S0(n1499) );
  HS65_GSS_XOR2X3 U1658 ( .A(n1500), .B(n1499), .Z(\mul_a2/fa1_s1[13] ) );
  HS65_GS_HA1X4 U1659 ( .A0(n1528), .B0(n1474), .CO(n1472), .S0(n1502) );
  HS65_GS_HA1X4 U1660 ( .A0(n1530), .B0(n1475), .CO(n1473), .S0(n1501) );
  HS65_GSS_XOR2X3 U1661 ( .A(n1502), .B(n1501), .Z(\mul_a2/fa1_s1[12] ) );
  HS65_GS_HA1X4 U1662 ( .A0(n1530), .B0(n1476), .CO(n1474), .S0(n1504) );
  HS65_GS_HA1X4 U1663 ( .A0(n1532), .B0(n1477), .CO(n1475), .S0(n1503) );
  HS65_GSS_XOR2X3 U1664 ( .A(n1504), .B(n1503), .Z(\mul_a2/fa1_s1[11] ) );
  HS65_GS_HA1X4 U1665 ( .A0(n1532), .B0(n1478), .CO(n1476), .S0(n1506) );
  HS65_GS_HA1X4 U1666 ( .A0(n1534), .B0(n1479), .CO(n1477), .S0(n1505) );
  HS65_GSS_XOR2X3 U1667 ( .A(n1506), .B(n1505), .Z(\mul_a2/fa1_s1[10] ) );
  HS65_GS_HA1X4 U1668 ( .A0(n1534), .B0(n1480), .CO(n1478), .S0(n1508) );
  HS65_GS_HA1X4 U1669 ( .A0(n1708), .B0(n1707), .CO(n1479), .S0(n1507) );
  HS65_GSS_XOR2X3 U1670 ( .A(n1508), .B(n1507), .Z(\mul_a2/fa1_s1[9] ) );
  HS65_GS_HA1X4 U1671 ( .A0(n1708), .B0(n1707), .CO(n1480), .S0(n1509) );
  HS65_GSS_XOR2X3 U1672 ( .A(n1509), .B(y_z2[0]), .Z(\mul_a2/fa1_s1[8] ) );
  HS65_GS_AND2X4 U1673 ( .A(n1482), .B(n1481), .Z(\mul_a2/fa1_c1[22] ) );
  HS65_GS_AND2X4 U1674 ( .A(n1484), .B(n1483), .Z(\mul_a2/fa1_c1[21] ) );
  HS65_GS_AND2X4 U1675 ( .A(n1486), .B(n1485), .Z(\mul_a2/fa1_c1[20] ) );
  HS65_GS_AND2X4 U1676 ( .A(n1488), .B(n1487), .Z(\mul_a2/fa1_c1[19] ) );
  HS65_GS_AND2X4 U1677 ( .A(n1490), .B(n1489), .Z(\mul_a2/fa1_c1[18] ) );
  HS65_GS_AND2X4 U1678 ( .A(n1492), .B(n1491), .Z(\mul_a2/fa1_c1[17] ) );
  HS65_GS_AND2X4 U1679 ( .A(n1494), .B(n1493), .Z(\mul_a2/fa1_c1[16] ) );
  HS65_GS_AND2X4 U1680 ( .A(n1496), .B(n1495), .Z(\mul_a2/fa1_c1[15] ) );
  HS65_GS_AND2X4 U1681 ( .A(n1498), .B(n1497), .Z(\mul_a2/fa1_c1[14] ) );
  HS65_GS_AND2X4 U1682 ( .A(n1500), .B(n1499), .Z(\mul_a2/fa1_c1[13] ) );
  HS65_GS_AND2X4 U1683 ( .A(n1502), .B(n1501), .Z(\mul_a2/fa1_c1[12] ) );
  HS65_GS_AND2X4 U1684 ( .A(n1504), .B(n1503), .Z(\mul_a2/fa1_c1[11] ) );
  HS65_GS_AND2X4 U1685 ( .A(n1506), .B(n1505), .Z(\mul_a2/fa1_c1[10] ) );
  HS65_GS_AND2X4 U1686 ( .A(n1508), .B(n1507), .Z(\mul_a2/fa1_c1[9] ) );
  HS65_GS_AND2X4 U1687 ( .A(n1509), .B(y_z2[0]), .Z(\mul_a2/fa1_c1[8] ) );
  HS65_GSS_XNOR2X3 U1688 ( .A(n1511), .B(n1510), .Z(\mul_a2/fa1_s2[28] ) );
  HS65_GSS_XNOR2X3 U1689 ( .A(n1513), .B(n1512), .Z(\mul_a2/fa1_s2[27] ) );
  HS65_GSS_XNOR2X3 U1690 ( .A(n1515), .B(n1514), .Z(\mul_a2/fa1_s2[26] ) );
  HS65_GSS_XNOR2X3 U1691 ( .A(n1517), .B(n1516), .Z(\mul_a2/fa1_s2[25] ) );
  HS65_GSS_XNOR2X3 U1692 ( .A(n1519), .B(n1518), .Z(\mul_a2/fa1_s2[24] ) );
  HS65_GSS_XNOR2X3 U1693 ( .A(n1521), .B(n1520), .Z(\mul_a2/fa1_s2[23] ) );
  HS65_GSS_XNOR2X3 U1694 ( .A(n1523), .B(n1522), .Z(\mul_a2/fa1_s2[22] ) );
  HS65_GSS_XNOR2X3 U1695 ( .A(n1525), .B(n1524), .Z(\mul_a2/fa1_s2[21] ) );
  HS65_GSS_XNOR2X3 U1696 ( .A(n1527), .B(n1526), .Z(\mul_a2/fa1_s2[20] ) );
  HS65_GSS_XNOR2X3 U1697 ( .A(n1529), .B(n1528), .Z(\mul_a2/fa1_s2[19] ) );
  HS65_GSS_XNOR2X3 U1698 ( .A(n1531), .B(n1530), .Z(\mul_a2/fa1_s2[18] ) );
  HS65_GSS_XNOR2X3 U1699 ( .A(n1533), .B(n1532), .Z(\mul_a2/fa1_s2[17] ) );
  HS65_GSS_XNOR2X3 U1700 ( .A(n1535), .B(n1534), .Z(\mul_a2/fa1_s2[16] ) );
  HS65_GSS_XNOR2X3 U1701 ( .A(n1536), .B(n1708), .Z(\mul_a2/fa1_s2[15] ) );
  HS65_GSS_XNOR2X3 U1702 ( .A(n1537), .B(n1707), .Z(\mul_a2/fa1_s2[14] ) );
  HS65_GS_FA1X4 U1703 ( .A0(n1540), .B0(n1539), .CI(n1538), .CO(n1549), .S0(
        n1560) );
  HS65_GS_FA1X4 U1704 ( .A0(n1543), .B0(n1542), .CI(n1541), .CO(n1553), .S0(
        n1544) );
  HS65_GS_IVX2 U1705 ( .A(n1544), .Z(n1558) );
  HS65_GS_FA1X4 U1706 ( .A0(n1547), .B0(n1546), .CI(n1545), .CO(n1542), .S0(
        n1557) );
  HS65_GS_FA1X4 U1707 ( .A0(n1550), .B0(n1549), .CI(n1548), .CO(n1546), .S0(
        n1556) );
  HS65_GS_FA1X4 U1708 ( .A0(n1553), .B0(n1552), .CI(n1551), .CO(n135), .S0(
        n1555) );
  HS65_GS_NAND3X2 U1709 ( .A(n1557), .B(n1556), .C(n1555), .Z(n1554) );
  HS65_GS_OAI12X3 U1710 ( .A(n1558), .B(n1554), .C(\mul_a2/result_sat[15] ), 
        .Z(n1617) );
  HS65_GS_NOR3X1 U1711 ( .A(n1557), .B(n1556), .C(n1555), .Z(n1559) );
  HS65_GS_AOI12X3 U1712 ( .A(n1559), .B(n1558), .C(\mul_a2/result_sat[15] ), 
        .Z(n1616) );
  HS65_GS_AO12X4 U1713 ( .A(n1560), .B(n1617), .C(n1616), .Z(
        \mul_a2/result_sat[14] ) );
  HS65_GS_FA1X4 U1714 ( .A0(n1563), .B0(n1562), .CI(n1561), .CO(n1539), .S0(
        n1564) );
  HS65_GS_AO12X4 U1715 ( .A(n1564), .B(n1617), .C(n1616), .Z(
        \mul_a2/result_sat[13] ) );
  HS65_GS_FA1X4 U1716 ( .A0(n1567), .B0(n1566), .CI(n1565), .CO(n1563), .S0(
        n1568) );
  HS65_GS_OA12X4 U1717 ( .A(n1616), .B(n1568), .C(n1617), .Z(
        \mul_a2/result_sat[12] ) );
  HS65_GS_FA1X4 U1718 ( .A0(n1571), .B0(n1570), .CI(n1569), .CO(n1567), .S0(
        n1572) );
  HS65_GS_OA12X4 U1719 ( .A(n1616), .B(n1572), .C(n1617), .Z(
        \mul_a2/result_sat[11] ) );
  HS65_GS_FA1X4 U1720 ( .A0(n1575), .B0(n1574), .CI(n1573), .CO(n1570), .S0(
        n1576) );
  HS65_GS_AO12X4 U1721 ( .A(n1576), .B(n1617), .C(n1616), .Z(
        \mul_a2/result_sat[10] ) );
  HS65_GS_FA1X4 U1722 ( .A0(n1579), .B0(n1578), .CI(n1577), .CO(n1575), .S0(
        n1580) );
  HS65_GS_AO12X4 U1723 ( .A(n1580), .B(n1617), .C(n1616), .Z(
        \mul_a2/result_sat[9] ) );
  HS65_GS_FA1X4 U1724 ( .A0(n1583), .B0(n1582), .CI(n1581), .CO(n1579), .S0(
        n1584) );
  HS65_GS_OA12X4 U1725 ( .A(n1616), .B(n1584), .C(n1617), .Z(
        \mul_a2/result_sat[8] ) );
  HS65_GS_FA1X4 U1726 ( .A0(n1587), .B0(n1586), .CI(n1585), .CO(n1583), .S0(
        n1588) );
  HS65_GS_OA12X4 U1727 ( .A(n1616), .B(n1588), .C(n1617), .Z(
        \mul_a2/result_sat[7] ) );
  HS65_GS_FA1X4 U1728 ( .A0(n1591), .B0(n1590), .CI(n1589), .CO(n1586), .S0(
        n1592) );
  HS65_GS_AO12X4 U1729 ( .A(n1592), .B(n1617), .C(n1616), .Z(
        \mul_a2/result_sat[6] ) );
  HS65_GS_FA1X4 U1730 ( .A0(n1595), .B0(n1594), .CI(n1593), .CO(n1590), .S0(
        n1596) );
  HS65_GS_AO12X4 U1731 ( .A(n1596), .B(n1617), .C(n1616), .Z(
        \mul_a2/result_sat[5] ) );
  HS65_GS_FA1X4 U1732 ( .A0(n1599), .B0(n1598), .CI(n1597), .CO(n1594), .S0(
        n1600) );
  HS65_GS_OA12X4 U1733 ( .A(n1616), .B(n1600), .C(n1617), .Z(
        \mul_a2/result_sat[4] ) );
  HS65_GS_FA1X4 U1734 ( .A0(n1603), .B0(n1602), .CI(n1601), .CO(n1598), .S0(
        n1604) );
  HS65_GS_AO12X4 U1735 ( .A(n1604), .B(n1617), .C(n1616), .Z(
        \mul_a2/result_sat[3] ) );
  HS65_GS_FA1X4 U1736 ( .A0(n1607), .B0(n1606), .CI(n1605), .CO(n1602), .S0(
        n1608) );
  HS65_GS_AO12X4 U1737 ( .A(n1608), .B(n1617), .C(n1616), .Z(
        \mul_a2/result_sat[2] ) );
  HS65_GS_FA1X4 U1738 ( .A0(n1611), .B0(n1610), .CI(n1609), .CO(n1606), .S0(
        n1612) );
  HS65_GS_AO12X4 U1739 ( .A(n1612), .B(n1617), .C(n1616), .Z(
        \mul_a2/result_sat[1] ) );
  HS65_GS_FA1X4 U1740 ( .A0(n1615), .B0(n1614), .CI(n1613), .CO(n1610), .S0(
        n1618) );
  HS65_GS_AO12X4 U1741 ( .A(n1618), .B(n1617), .C(n1616), .Z(
        \mul_a2/result_sat[0] ) );
  HS65_GSS_XNOR2X3 U1742 ( .A(n1619), .B(n1639), .Z(\mul_a1/fa1_s0[16] ) );
  HS65_GSS_XNOR2X3 U1743 ( .A(n1620), .B(n1641), .Z(\mul_a1/fa1_s0[15] ) );
  HS65_GSS_XNOR2X3 U1744 ( .A(n1621), .B(n1643), .Z(\mul_a1/fa1_s0[14] ) );
  HS65_GSS_XNOR2X3 U1745 ( .A(n1622), .B(n1645), .Z(\mul_a1/fa1_s0[13] ) );
  HS65_GSS_XNOR2X3 U1746 ( .A(n1623), .B(n1647), .Z(\mul_a1/fa1_s0[12] ) );
  HS65_GSS_XNOR2X3 U1747 ( .A(n1624), .B(n1649), .Z(\mul_a1/fa1_s0[11] ) );
  HS65_GSS_XNOR2X3 U1748 ( .A(n1625), .B(n1651), .Z(\mul_a1/fa1_s0[10] ) );
  HS65_GSS_XNOR2X3 U1749 ( .A(n1626), .B(n1653), .Z(\mul_a1/fa1_s0[9] ) );
  HS65_GSS_XNOR2X3 U1750 ( .A(n1627), .B(n1655), .Z(\mul_a1/fa1_s0[8] ) );
  HS65_GSS_XNOR2X3 U1751 ( .A(n1628), .B(n1657), .Z(\mul_a1/fa1_s0[7] ) );
  HS65_GSS_XNOR2X3 U1752 ( .A(n1629), .B(n1659), .Z(\mul_a1/fa1_s0[6] ) );
  HS65_GSS_XNOR2X3 U1753 ( .A(n1630), .B(n1661), .Z(\mul_a1/fa1_s0[5] ) );
  HS65_GSS_XNOR2X3 U1754 ( .A(n1631), .B(n1713), .Z(\mul_a1/fa1_s0[4] ) );
  HS65_GS_AND2X4 U1755 ( .A(n1632), .B(y_z1[14]), .Z(\mul_a1/fa1_c0[17] ) );
  HS65_GSS_XNOR2X3 U1756 ( .A(y_z1[15]), .B(n1633), .Z(\C55/DATA4_28 ) );
  HS65_GS_HA1X4 U1757 ( .A0(n1635), .B0(n1634), .CO(n1633), .S0(\C55/DATA4_27 ) );
  HS65_GS_HA1X4 U1758 ( .A0(n1637), .B0(n1636), .CO(n1634), .S0(\C55/DATA4_26 ) );
  HS65_GS_HA1X4 U1759 ( .A0(n1639), .B0(n1638), .CO(n1636), .S0(\C55/DATA4_25 ) );
  HS65_GS_HA1X4 U1760 ( .A0(n1641), .B0(n1640), .CO(n1638), .S0(\C55/DATA4_24 ) );
  HS65_GS_HA1X4 U1761 ( .A0(n1643), .B0(n1642), .CO(n1640), .S0(\C55/DATA4_23 ) );
  HS65_GS_HA1X4 U1762 ( .A0(n1645), .B0(n1644), .CO(n1642), .S0(\C55/DATA4_22 ) );
  HS65_GS_HA1X4 U1763 ( .A0(n1647), .B0(n1646), .CO(n1644), .S0(\C55/DATA4_21 ) );
  HS65_GS_HA1X4 U1764 ( .A0(n1649), .B0(n1648), .CO(n1646), .S0(\C55/DATA4_20 ) );
  HS65_GS_HA1X4 U1765 ( .A0(n1651), .B0(n1650), .CO(n1648), .S0(\C55/DATA4_19 ) );
  HS65_GS_HA1X4 U1766 ( .A0(n1653), .B0(n1652), .CO(n1650), .S0(\C55/DATA4_18 ) );
  HS65_GS_HA1X4 U1767 ( .A0(n1655), .B0(n1654), .CO(n1652), .S0(\C55/DATA4_17 ) );
  HS65_GS_HA1X4 U1768 ( .A0(n1657), .B0(n1656), .CO(n1654), .S0(\C55/DATA4_16 ) );
  HS65_GS_HA1X4 U1769 ( .A0(n1659), .B0(n1658), .CO(n1656), .S0(\C55/DATA4_15 ) );
  HS65_GS_HA1X4 U1770 ( .A0(n1661), .B0(n1660), .CO(n1658), .S0(\C55/DATA4_14 ) );
  HS65_GS_HA1X4 U1771 ( .A0(n1713), .B0(n1712), .CO(n1660), .S0(\C55/DATA4_13 ) );
  HS65_GSS_XNOR2X3 U1772 ( .A(x_reg2[15]), .B(n1662), .Z(\C43/DATA4_22 ) );
  HS65_GS_HA1X4 U1773 ( .A0(n1727), .B0(n1663), .CO(n1662), .S0(\C43/DATA4_21 ) );
  HS65_GS_HA1X4 U1774 ( .A0(n1728), .B0(n1664), .CO(n1663), .S0(\C43/DATA4_20 ) );
  HS65_GS_HA1X4 U1775 ( .A0(n1726), .B0(n1665), .CO(n1664), .S0(\C43/DATA4_19 ) );
  HS65_GS_HA1X4 U1776 ( .A0(n1725), .B0(n1666), .CO(n1665), .S0(\C43/DATA4_18 ) );
  HS65_GS_HA1X4 U1777 ( .A0(n1724), .B0(n1667), .CO(n1666), .S0(\C43/DATA4_17 ) );
  HS65_GS_HA1X4 U1778 ( .A0(n1723), .B0(n1668), .CO(n1667), .S0(\C43/DATA4_16 ) );
  HS65_GS_HA1X4 U1779 ( .A0(n1722), .B0(n1669), .CO(n1668), .S0(\C43/DATA4_15 ) );
  HS65_GS_HA1X4 U1780 ( .A0(n1721), .B0(n1670), .CO(n1669), .S0(\C43/DATA4_14 ) );
  HS65_GS_HA1X4 U1781 ( .A0(n1720), .B0(n1671), .CO(n1670), .S0(\C43/DATA4_13 ) );
  HS65_GS_HA1X4 U1782 ( .A0(n1719), .B0(n1672), .CO(n1671), .S0(\C43/DATA4_12 ) );
  HS65_GS_HA1X4 U1783 ( .A0(n1718), .B0(n1673), .CO(n1672), .S0(\C43/DATA4_11 ) );
  HS65_GS_HA1X4 U1784 ( .A0(n1717), .B0(n1674), .CO(n1673), .S0(\C43/DATA4_10 ) );
  HS65_GS_HA1X4 U1785 ( .A0(n1716), .B0(n1675), .CO(n1674), .S0(\C43/DATA4_9 )
         );
  HS65_GS_HA1X4 U1786 ( .A0(n1715), .B0(n1676), .CO(n1675), .S0(\C43/DATA4_8 )
         );
  HS65_GS_HA1X4 U1787 ( .A0(n1714), .B0(n1677), .CO(n1676), .S0(
        \mul_b2/fa1_s1[7] ) );
  HS65_GSS_XNOR2X3 U1788 ( .A(x_z2[15]), .B(n1678), .Z(\C33/DATA4_20 ) );
  HS65_GS_HA1X4 U1789 ( .A0(n1680), .B0(n1679), .CO(n1678), .S0(\C33/DATA4_19 ) );
  HS65_GS_HA1X4 U1790 ( .A0(n1682), .B0(n1681), .CO(n1679), .S0(\C33/DATA4_18 ) );
  HS65_GS_HA1X4 U1791 ( .A0(n1684), .B0(n1683), .CO(n1681), .S0(\C33/DATA4_17 ) );
  HS65_GS_HA1X4 U1792 ( .A0(n1686), .B0(n1685), .CO(n1683), .S0(\C33/DATA4_16 ) );
  HS65_GS_HA1X4 U1793 ( .A0(n1688), .B0(n1687), .CO(n1685), .S0(\C33/DATA4_15 ) );
  HS65_GS_HA1X4 U1794 ( .A0(n1690), .B0(n1689), .CO(n1687), .S0(\C33/DATA4_14 ) );
  HS65_GS_HA1X4 U1795 ( .A0(n1692), .B0(n1691), .CO(n1689), .S0(\C33/DATA4_13 ) );
  HS65_GS_HA1X4 U1796 ( .A0(n1694), .B0(n1693), .CO(n1691), .S0(\C33/DATA4_12 ) );
  HS65_GS_HA1X4 U1797 ( .A0(n1696), .B0(n1695), .CO(n1693), .S0(\C33/DATA4_11 ) );
  HS65_GS_HA1X4 U1798 ( .A0(n1698), .B0(n1697), .CO(n1695), .S0(\C33/DATA4_10 ) );
  HS65_GS_HA1X4 U1799 ( .A0(n1700), .B0(n1699), .CO(n1697), .S0(\C33/DATA4_9 )
         );
  HS65_GS_HA1X4 U1800 ( .A0(n1702), .B0(n1701), .CO(n1699), .S0(\C33/DATA4_8 )
         );
  HS65_GS_HA1X4 U1801 ( .A0(n1704), .B0(n1703), .CO(n1701), .S0(\C33/DATA4_7 )
         );
  HS65_GS_HA1X4 U1802 ( .A0(n1706), .B0(n1705), .CO(n1703), .S0(\C33/DATA4_6 )
         );
  HS65_GS_HA1X4 U1803 ( .A0(n1708), .B0(n1707), .CO(n1381), .S0(\C64/DATA4_13 ) );
  HS65_GS_HA1X4 U1804 ( .A0(n1710), .B0(n1709), .CO(n1711), .S0(n981) );
  HS65_GSS_XNOR2X3 U1805 ( .A(y_z2[15]), .B(n1711), .Z(\mul_a2/fa1_c1[24] ) );
  HS65_GS_HA1X4 U1806 ( .A0(n1713), .B0(n1712), .CO(n1415), .S0(\C53/DATA4_10 ) );
  HS65_GS_HA1X4 U1807 ( .A0(n1349), .B0(n1347), .CO(n1005), .S0(
        \mul_b1/fa1_s1[7] ) );
  HS65_GS_AOI12X2 U1808 ( .A(n1714), .B(n1716), .C(\mul_b2/fa1_c0[5] ), .Z(
        \mul_b2/fa1_s0[5] ) );
  HS65_GS_AOI12X2 U1809 ( .A(n1715), .B(n1717), .C(\mul_b2/fa1_c0[6] ), .Z(
        \mul_b2/fa1_s0[6] ) );
  HS65_GS_AOI12X2 U1810 ( .A(n1716), .B(n1718), .C(\mul_b2/fa1_c0[7] ), .Z(
        \mul_b2/fa1_s0[7] ) );
  HS65_GS_AOI12X2 U1811 ( .A(n1717), .B(n1719), .C(\mul_b2/fa1_c0[8] ), .Z(
        \mul_b2/fa1_s0[8] ) );
  HS65_GS_AOI12X2 U1812 ( .A(n1718), .B(n1720), .C(\mul_b2/fa1_c0[9] ), .Z(
        \mul_b2/fa1_s0[9] ) );
  HS65_GS_AOI12X2 U1813 ( .A(n1719), .B(n1721), .C(\mul_b2/fa1_c0[10] ), .Z(
        \mul_b2/fa1_s0[10] ) );
  HS65_GS_AOI12X2 U1814 ( .A(n1720), .B(n1722), .C(\mul_b2/fa1_c0[11] ), .Z(
        \mul_b2/fa1_s0[11] ) );
  HS65_GS_AOI12X2 U1815 ( .A(n1721), .B(n1723), .C(\mul_b2/fa1_c0[12] ), .Z(
        \mul_b2/fa1_s0[12] ) );
  HS65_GS_AOI12X2 U1816 ( .A(n1722), .B(n1724), .C(\mul_b2/fa1_c0[13] ), .Z(
        \mul_b2/fa1_s0[13] ) );
  HS65_GS_AOI12X2 U1817 ( .A(n1723), .B(n1725), .C(\mul_b2/fa1_c0[14] ), .Z(
        \mul_b2/fa1_s0[14] ) );
  HS65_GS_AOI12X2 U1818 ( .A(n1724), .B(n1726), .C(\mul_b2/fa1_c0[15] ), .Z(
        \mul_b2/fa1_s0[15] ) );
  HS65_GS_AOI12X2 U1819 ( .A(n1725), .B(n1728), .C(\mul_b2/fa1_c0[16] ), .Z(
        \mul_b2/fa1_s0[16] ) );
  HS65_GS_AOI12X2 U1820 ( .A(n1726), .B(n1727), .C(\mul_b2/fa1_c0[17] ), .Z(
        \mul_b2/fa1_s0[17] ) );
  HS65_GS_AOI12X2 U1821 ( .A(n1728), .B(n1727), .C(\mul_b2/fa1_c0[18] ), .Z(
        \mul_b2/fa1_s0[18] ) );
  HS65_GS_AOI12X2 U1822 ( .A(n1731), .B(n1730), .C(n1729), .Z(n1732) );
  HS65_GS_AOI12X2 U1823 ( .A(n1732), .B(n1745), .C(n1744), .Z(
        \mul_a1/result_sat[0] ) );
  HS65_GS_OAI112X1 U1824 ( .A(n1735), .B(n1734), .C(n1745), .D(n1733), .Z(
        n1736) );
  HS65_GS_NOR2AX3 U1825 ( .A(n1736), .B(n1744), .Z(\mul_a1/result_sat[3] ) );
  HS65_GS_OAI112X1 U1826 ( .A(n1739), .B(n1738), .C(n1745), .D(n1737), .Z(
        n1740) );
  HS65_GS_NOR2AX3 U1827 ( .A(n1740), .B(n1744), .Z(\mul_a1/result_sat[6] ) );
  HS65_GS_AOI12X2 U1828 ( .A(n1743), .B(n1742), .C(n1741), .Z(n1746) );
  HS65_GS_AOI12X2 U1829 ( .A(n1746), .B(n1745), .C(n1744), .Z(
        \mul_a1/result_sat[12] ) );
  HS65_GS_AOI12X2 U1830 ( .A(n1749), .B(n1748), .C(n1747), .Z(n1751) );
  HS65_GS_IVX2 U1831 ( .A(n1750), .Z(n1779) );
  HS65_GS_AOI12X2 U1832 ( .A(n1751), .B(n1780), .C(n1779), .Z(
        \mul_b1/result_sat[0] ) );
  HS65_GS_AOI12X2 U1833 ( .A(n1754), .B(n1753), .C(n1752), .Z(n1755) );
  HS65_GS_AOI12X2 U1834 ( .A(n1755), .B(n1780), .C(n1779), .Z(
        \mul_b1/result_sat[1] ) );
  HS65_GS_AOI12X2 U1835 ( .A(n1758), .B(n1757), .C(n1756), .Z(n1759) );
  HS65_GS_AOI12X2 U1836 ( .A(n1759), .B(n1780), .C(n1779), .Z(
        \mul_b1/result_sat[2] ) );
  HS65_GS_AOI12X2 U1837 ( .A(n1762), .B(n1761), .C(n1760), .Z(n1763) );
  HS65_GS_AOI12X2 U1838 ( .A(n1763), .B(n1780), .C(n1779), .Z(
        \mul_b1/result_sat[3] ) );
  HS65_GS_AOI12X2 U1839 ( .A(n1766), .B(n1765), .C(n1764), .Z(n1767) );
  HS65_GS_AOI12X2 U1840 ( .A(n1767), .B(n1780), .C(n1779), .Z(
        \mul_b1/result_sat[4] ) );
  HS65_GS_AOI12X2 U1841 ( .A(n1770), .B(n1769), .C(n1768), .Z(n1771) );
  HS65_GS_AOI12X2 U1842 ( .A(n1771), .B(n1780), .C(n1779), .Z(
        \mul_b1/result_sat[5] ) );
  HS65_GS_AOI12X2 U1843 ( .A(n1774), .B(n1773), .C(n1772), .Z(n1775) );
  HS65_GS_AOI12X2 U1844 ( .A(n1775), .B(n1780), .C(n1779), .Z(
        \mul_b1/result_sat[6] ) );
  HS65_GS_AOI12X2 U1845 ( .A(n1778), .B(n1777), .C(n1776), .Z(n1781) );
  HS65_GS_AOI12X2 U1846 ( .A(n1781), .B(n1780), .C(n1779), .Z(
        \mul_b1/result_sat[7] ) );
  HS65_GS_AOI12X2 U1847 ( .A(n1784), .B(n1783), .C(n1782), .Z(n1841) );
endmodule


module opti_sos_1 ( clk, rst_n, data_in, valid_in, b0, b1, b2, a1, a2, 
        data_out, valid_out );
  input [15:0] data_in;
  input [15:0] b0;
  input [15:0] b1;
  input [15:0] b2;
  input [15:0] a1;
  input [15:0] a2;
  output [15:0] data_out;
  input clk, rst_n, valid_in;
  output valid_out;
  wire   valid_T1, valid_T3, valid_T2, \mul_b0/result_sat[15] ,
         \mul_b0/result_sat[14] , \mul_b0/result_sat[13] ,
         \mul_b0/result_sat[12] , \mul_b0/result_sat[11] ,
         \mul_b0/result_sat[10] , \mul_b0/result_sat[9] ,
         \mul_b0/result_sat[8] , \mul_b0/result_sat[7] ,
         \mul_b0/result_sat[6] , \mul_b0/result_sat[5] ,
         \mul_b0/result_sat[4] , \mul_b0/result_sat[3] ,
         \mul_b0/result_sat[2] , \mul_b0/result_sat[1] ,
         \mul_b0/result_sat[0] , \mul_b0/fa1_s2_r[33] , \mul_b0/fa1_s2_r[32] ,
         \mul_b0/fa1_s2_r[31] , \mul_b0/fa1_s2_r[30] , \mul_b0/fa1_s2_r[29] ,
         \mul_b0/fa1_s2_r[28] , \mul_b0/fa1_s2_r[27] , \mul_b0/fa1_s2_r[26] ,
         \mul_b0/fa1_s2_r[25] , \mul_b0/fa1_s2_r[24] , \mul_b0/fa1_s2_r[23] ,
         \mul_b0/fa1_s2_r[22] , \mul_b0/fa1_s2_r[21] , \mul_b0/fa1_s2_r[20] ,
         \mul_b0/fa1_s2_r[19] , \mul_b0/fa1_s2_r[18] , \mul_b0/fa1_s2_r[17] ,
         \mul_b0/fa1_s2_r[16] , \mul_b0/fa1_s2_r[15] , \mul_b0/fa1_s2_r[14] ,
         \mul_b0/fa1_s2_r[13] , \mul_b0/fa1_s2_r[12] , \mul_b0/fa1_s1_r[33] ,
         \mul_b0/fa1_s1_r[32] , \mul_b0/fa1_s1_r[31] , \mul_b0/fa1_s1_r[30] ,
         \mul_b0/fa1_s1_r[29] , \mul_b0/fa1_s1_r[28] , \mul_b0/fa1_s1_r[27] ,
         \mul_b0/fa1_s1_r[26] , \mul_b0/fa1_s1_r[25] , \mul_b0/fa1_s1_r[24] ,
         \mul_b0/fa1_s1_r[23] , \mul_b0/fa1_s1_r[22] , \mul_b0/fa1_s1_r[21] ,
         \mul_b0/fa1_s1_r[20] , \mul_b0/fa1_s1_r[19] , \mul_b0/fa1_s1_r[18] ,
         \mul_b0/fa1_s1_r[17] , \mul_b0/fa1_s1_r[16] , \mul_b0/fa1_s1_r[15] ,
         \mul_b0/fa1_s1_r[14] , \mul_b0/fa1_s1_r[13] , \mul_b0/fa1_s1_r[12] ,
         \mul_b0/fa1_s1_r[11] , \mul_b0/fa1_s1_r[10] , \mul_b0/fa1_s1_r[9] ,
         \mul_b0/fa1_s1_r[8] , \mul_b0/fa1_c0_r[20] , \mul_b0/fa1_c0_r[19] ,
         \mul_b0/fa1_c0_r[18] , \mul_b0/fa1_c0_r[17] , \mul_b0/fa1_c0_r[16] ,
         \mul_b0/fa1_c0_r[15] , \mul_b0/fa1_c0_r[14] , \mul_b0/fa1_c0_r[13] ,
         \mul_b0/fa1_c0_r[12] , \mul_b0/fa1_c0_r[11] , \mul_b0/fa1_c0_r[10] ,
         \mul_b0/fa1_c0_r[9] , \mul_b0/fa1_c0_r[8] , \mul_b0/fa1_c0_r[7] ,
         \mul_b0/fa1_c0_r[6] , \mul_b0/fa1_c0_r[5] , \mul_b0/fa1_s0_r[33] ,
         \mul_b0/fa1_s0_r[32] , \mul_b0/fa1_s0_r[31] , \mul_b0/fa1_s0_r[30] ,
         \mul_b0/fa1_s0_r[29] , \mul_b0/fa1_s0_r[28] , \mul_b0/fa1_s0_r[27] ,
         \mul_b0/fa1_s0_r[26] , \mul_b0/fa1_s0_r[25] , \mul_b0/fa1_s0_r[24] ,
         \mul_b0/fa1_s0_r[23] , \mul_b0/fa1_s0_r[22] , \mul_b0/fa1_s0_r[21] ,
         \mul_b0/fa1_s0_r[20] , \mul_b0/fa1_s0_r[19] , \mul_b0/fa1_s0_r[18] ,
         \mul_b0/fa1_s0_r[17] , \mul_b0/fa1_s0_r[16] , \mul_b0/fa1_s0_r[15] ,
         \mul_b0/fa1_s0_r[14] , \mul_b0/fa1_s0_r[13] , \mul_b0/fa1_s0_r[12] ,
         \mul_b0/fa1_s0_r[11] , \mul_b0/fa1_s0_r[10] , \mul_b0/fa1_s0_r[9] ,
         \mul_b0/fa1_s0_r[8] , \mul_b0/fa1_s0_r[7] , \mul_b0/fa1_s0_r[6] ,
         \mul_b0/fa1_c0[20] , \mul_b0/fa1_c0[19] , \mul_b0/fa1_c0[18] ,
         \mul_b0/fa1_c0[17] , \mul_b0/fa1_c0[16] , \mul_b0/fa1_c0[15] ,
         \mul_b0/fa1_c0[14] , \mul_b0/fa1_c0[13] , \mul_b0/fa1_c0[12] ,
         \mul_b0/fa1_c0[11] , \mul_b0/fa1_c0[10] , \mul_b0/fa1_c0[9] ,
         \mul_b0/fa1_c0[8] , \mul_b0/fa1_c0[7] , \mul_b0/fa1_c0[6] ,
         \mul_b0/fa1_c0[5] , \mul_b0/fa1_s0[31] , \mul_b0/fa1_s0[20] ,
         \mul_b0/fa1_s0[19] , \mul_b0/fa1_s0[18] , \mul_b0/fa1_s0[17] ,
         \mul_b0/fa1_s0[16] , \mul_b0/fa1_s0[15] , \mul_b0/fa1_s0[14] ,
         \mul_b0/fa1_s0[13] , \mul_b0/fa1_s0[12] , \mul_b0/fa1_s0[11] ,
         \mul_b0/fa1_s0[10] , \mul_b0/fa1_s0[9] , \mul_b0/fa1_s0[8] ,
         \mul_b0/fa1_s0[7] , \mul_b0/fa1_s0[6] , \mul_b1/result_sat[15] ,
         \mul_b1/result_sat[14] , \mul_b1/result_sat[13] ,
         \mul_b1/result_sat[12] , \mul_b1/result_sat[11] ,
         \mul_b1/result_sat[10] , \mul_b1/result_sat[9] ,
         \mul_b1/result_sat[8] , \mul_b1/result_sat[7] ,
         \mul_b1/result_sat[6] , \mul_b1/result_sat[5] ,
         \mul_b1/result_sat[4] , \mul_b1/result_sat[3] ,
         \mul_b1/result_sat[2] , \mul_b1/result_sat[1] ,
         \mul_b1/result_sat[0] , \mul_b1/fa1_c2_r[28] , \mul_b1/fa1_c2_r[27] ,
         \mul_b1/fa1_c2_r[26] , \mul_b1/fa1_c2_r[25] , \mul_b1/fa1_c2_r[24] ,
         \mul_b1/fa1_c2_r[23] , \mul_b1/fa1_c2_r[22] , \mul_b1/fa1_c2_r[21] ,
         \mul_b1/fa1_c2_r[20] , \mul_b1/fa1_c2_r[19] , \mul_b1/fa1_c2_r[18] ,
         \mul_b1/fa1_c2_r[17] , \mul_b1/fa1_c2_r[16] , \mul_b1/fa1_c2_r[15] ,
         \mul_b1/fa1_c2_r[14] , \mul_b1/fa1_s2_r[33] , \mul_b1/fa1_s2_r[32] ,
         \mul_b1/fa1_s2_r[31] , \mul_b1/fa1_s2_r[30] , \mul_b1/fa1_s2_r[29] ,
         \mul_b1/fa1_s2_r[28] , \mul_b1/fa1_s2_r[27] , \mul_b1/fa1_s2_r[26] ,
         \mul_b1/fa1_s2_r[25] , \mul_b1/fa1_s2_r[24] , \mul_b1/fa1_s2_r[23] ,
         \mul_b1/fa1_s2_r[22] , \mul_b1/fa1_s2_r[21] , \mul_b1/fa1_s2_r[20] ,
         \mul_b1/fa1_s2_r[19] , \mul_b1/fa1_s2_r[18] , \mul_b1/fa1_s2_r[17] ,
         \mul_b1/fa1_s2_r[16] , \mul_b1/fa1_s2_r[15] , \mul_b1/fa1_s2_r[14] ,
         \mul_b1/fa1_s2_r[13] , \mul_b1/fa1_c1_r[32] , \mul_b1/fa1_c1_r[31] ,
         \mul_b1/fa1_c1_r[30] , \mul_b1/fa1_c1_r[29] , \mul_b1/fa1_c1_r[28] ,
         \mul_b1/fa1_c1_r[27] , \mul_b1/fa1_c1_r[26] , \mul_b1/fa1_c1_r[25] ,
         \mul_b1/fa1_c1_r[24] , \mul_b1/fa1_c1_r[23] , \mul_b1/fa1_c1_r[22] ,
         \mul_b1/fa1_c1_r[21] , \mul_b1/fa1_c1_r[20] , \mul_b1/fa1_c1_r[19] ,
         \mul_b1/fa1_c1_r[18] , \mul_b1/fa1_c1_r[17] , \mul_b1/fa1_c1_r[16] ,
         \mul_b1/fa1_c1_r[15] , \mul_b1/fa1_c1_r[14] , \mul_b1/fa1_c1_r[13] ,
         \mul_b1/fa1_c1_r[12] , \mul_b1/fa1_c1_r[11] , \mul_b1/fa1_c1_r[10] ,
         \mul_b1/fa1_c1_r[9] , \mul_b1/fa1_c1_r[8] , \mul_b1/fa1_s1_r[22] ,
         \mul_b1/fa1_s1_r[21] , \mul_b1/fa1_s1_r[20] , \mul_b1/fa1_s1_r[19] ,
         \mul_b1/fa1_s1_r[18] , \mul_b1/fa1_s1_r[17] , \mul_b1/fa1_s1_r[16] ,
         \mul_b1/fa1_s1_r[15] , \mul_b1/fa1_s1_r[14] , \mul_b1/fa1_s1_r[13] ,
         \mul_b1/fa1_s1_r[12] , \mul_b1/fa1_s1_r[11] , \mul_b1/fa1_s1_r[10] ,
         \mul_b1/fa1_s1_r[9] , \mul_b1/fa1_s1_r[8] , \mul_b1/fa1_s1_r[7] ,
         \mul_b1/fa1_s1_r[6] , \mul_b1/fa1_c0_r[32] , \mul_b1/fa1_c0_r[31] ,
         \mul_b1/fa1_c0_r[30] , \mul_b1/fa1_c0_r[29] , \mul_b1/fa1_c0_r[28] ,
         \mul_b1/fa1_c0_r[27] , \mul_b1/fa1_c0_r[26] , \mul_b1/fa1_c0_r[25] ,
         \mul_b1/fa1_c0_r[24] , \mul_b1/fa1_c0_r[23] , \mul_b1/fa1_c0_r[22] ,
         \mul_b1/fa1_c0_r[21] , \mul_b1/fa1_c0_r[20] , \mul_b1/fa1_c0_r[19] ,
         \mul_b1/fa1_c0_r[18] , \mul_b1/fa1_c0_r[17] , \mul_b1/fa1_c0_r[16] ,
         \mul_b1/fa1_c0_r[15] , \mul_b1/fa1_c0_r[14] , \mul_b1/fa1_c0_r[13] ,
         \mul_b1/fa1_c0_r[12] , \mul_b1/fa1_c0_r[11] , \mul_b1/fa1_c0_r[10] ,
         \mul_b1/fa1_c0_r[9] , \mul_b1/fa1_c0_r[8] , \mul_b1/fa1_c0_r[7] ,
         \mul_b1/fa1_c0_r[6] , \mul_b1/fa1_c0_r[5] , \mul_b1/fa1_c0_r[4] ,
         \mul_b1/fa1_c0_r[3] , \mul_b1/fa1_c0_r[2] , \mul_b1/fa1_s0_r[33] ,
         \mul_b1/fa1_s0_r[32] , \mul_b1/fa1_s0_r[31] , \mul_b1/fa1_s0_r[30] ,
         \mul_b1/fa1_s0_r[29] , \mul_b1/fa1_s0_r[28] , \mul_b1/fa1_s0_r[27] ,
         \mul_b1/fa1_s0_r[26] , \mul_b1/fa1_s0_r[25] , \mul_b1/fa1_s0_r[24] ,
         \mul_b1/fa1_s0_r[23] , \mul_b1/fa1_s0_r[22] , \mul_b1/fa1_s0_r[21] ,
         \mul_b1/fa1_s0_r[20] , \mul_b1/fa1_s0_r[19] , \mul_b1/fa1_s0_r[18] ,
         \mul_b1/fa1_s0_r[17] , \mul_b1/fa1_s0_r[16] , \mul_b1/fa1_s0_r[15] ,
         \mul_b1/fa1_s0_r[14] , \mul_b1/fa1_s0_r[13] , \mul_b1/fa1_s0_r[12] ,
         \mul_b1/fa1_s0_r[11] , \mul_b1/fa1_s0_r[10] , \mul_b1/fa1_s0_r[9] ,
         \mul_b1/fa1_s0_r[8] , \mul_b1/fa1_s0_r[7] , \mul_b1/fa1_s0_r[6] ,
         \mul_b1/fa1_s0_r[5] , \mul_b1/fa1_s0_r[4] , \mul_b1/fa1_s0_r[3] ,
         \mul_b1/fa1_c2[28] , \mul_b1/fa1_c2[27] , \mul_b1/fa1_c2[26] ,
         \mul_b1/fa1_c2[25] , \mul_b1/fa1_c2[24] , \mul_b1/fa1_c2[23] ,
         \mul_b1/fa1_c2[22] , \mul_b1/fa1_c2[21] , \mul_b1/fa1_c2[20] ,
         \mul_b1/fa1_c2[19] , \mul_b1/fa1_c2[18] , \mul_b1/fa1_c2[17] ,
         \mul_b1/fa1_c2[16] , \mul_b1/fa1_c2[15] , \mul_b1/fa1_c2[14] ,
         \mul_b1/fa1_s2[29] , \mul_b1/fa1_s2[28] , \mul_b1/fa1_s2[27] ,
         \mul_b1/fa1_s2[26] , \mul_b1/fa1_s2[25] , \mul_b1/fa1_s2[24] ,
         \mul_b1/fa1_s2[23] , \mul_b1/fa1_s2[22] , \mul_b1/fa1_s2[21] ,
         \mul_b1/fa1_s2[20] , \mul_b1/fa1_s2[19] , \mul_b1/fa1_s2[18] ,
         \mul_b1/fa1_s2[17] , \mul_b1/fa1_s2[16] , \mul_b1/fa1_s2[15] ,
         \mul_b1/fa1_s2[14] , \mul_b1/fa1_c1[22] , \mul_b1/fa1_c1[21] ,
         \mul_b1/fa1_c1[20] , \mul_b1/fa1_c1[19] , \mul_b1/fa1_c1[18] ,
         \mul_b1/fa1_c1[17] , \mul_b1/fa1_c1[16] , \mul_b1/fa1_c1[15] ,
         \mul_b1/fa1_c1[14] , \mul_b1/fa1_c1[13] , \mul_b1/fa1_c1[12] ,
         \mul_b1/fa1_c1[11] , \mul_b1/fa1_c1[10] , \mul_b1/fa1_c1[9] ,
         \mul_b1/fa1_c1[8] , \mul_b1/fa1_s1[22] , \mul_b1/fa1_s1[21] ,
         \mul_b1/fa1_s1[20] , \mul_b1/fa1_s1[19] , \mul_b1/fa1_s1[18] ,
         \mul_b1/fa1_s1[17] , \mul_b1/fa1_s1[16] , \mul_b1/fa1_s1[15] ,
         \mul_b1/fa1_s1[14] , \mul_b1/fa1_s1[13] , \mul_b1/fa1_s1[12] ,
         \mul_b1/fa1_s1[11] , \mul_b1/fa1_s1[10] , \mul_b1/fa1_s1[9] ,
         \mul_b1/fa1_s1[8] , \mul_b1/fa1_c0[18] , \mul_b1/fa1_c0[17] ,
         \mul_b1/fa1_c0[16] , \mul_b1/fa1_c0[15] , \mul_b1/fa1_c0[14] ,
         \mul_b1/fa1_c0[13] , \mul_b1/fa1_c0[12] , \mul_b1/fa1_c0[11] ,
         \mul_b1/fa1_c0[10] , \mul_b1/fa1_c0[9] , \mul_b1/fa1_c0[8] ,
         \mul_b1/fa1_c0[7] , \mul_b1/fa1_c0[6] , \mul_b1/fa1_c0[5] ,
         \mul_b1/fa1_c0[4] , \mul_b1/fa1_s0[28] , \mul_b1/fa1_s0[20] ,
         \mul_b1/fa1_s0[19] , \mul_b1/fa1_s0[18] , \mul_b1/fa1_s0[17] ,
         \mul_b1/fa1_s0[16] , \mul_b1/fa1_s0[15] , \mul_b1/fa1_s0[14] ,
         \mul_b1/fa1_s0[13] , \mul_b1/fa1_s0[12] , \mul_b1/fa1_s0[11] ,
         \mul_b1/fa1_s0[10] , \mul_b1/fa1_s0[9] , \mul_b1/fa1_s0[8] ,
         \mul_b1/fa1_s0[7] , \mul_b1/fa1_s0[6] , \mul_b1/fa1_s0[5] ,
         \mul_b1/fa1_s0[4] , \mul_b1/fa1_s0[3] , \mul_b1/fa1_s0[1] ,
         \mul_b1/fa1_s0[0] , \mul_b2/result_sat[15] , \mul_b2/result_sat[14] ,
         \mul_b2/result_sat[13] , \mul_b2/result_sat[12] ,
         \mul_b2/result_sat[11] , \mul_b2/result_sat[10] ,
         \mul_b2/result_sat[9] , \mul_b2/result_sat[8] ,
         \mul_b2/result_sat[7] , \mul_b2/result_sat[6] ,
         \mul_b2/result_sat[5] , \mul_b2/result_sat[4] ,
         \mul_b2/result_sat[3] , \mul_b2/result_sat[2] ,
         \mul_b2/result_sat[1] , \mul_b2/result_sat[0] , \mul_b2/fa1_s2_r[33] ,
         \mul_b2/fa1_s2_r[32] , \mul_b2/fa1_s2_r[31] , \mul_b2/fa1_s2_r[30] ,
         \mul_b2/fa1_s2_r[29] , \mul_b2/fa1_s2_r[28] , \mul_b2/fa1_s2_r[27] ,
         \mul_b2/fa1_s2_r[26] , \mul_b2/fa1_s2_r[25] , \mul_b2/fa1_s2_r[24] ,
         \mul_b2/fa1_s2_r[23] , \mul_b2/fa1_s2_r[22] , \mul_b2/fa1_s2_r[21] ,
         \mul_b2/fa1_s2_r[20] , \mul_b2/fa1_s2_r[19] , \mul_b2/fa1_s2_r[18] ,
         \mul_b2/fa1_s2_r[17] , \mul_b2/fa1_s2_r[16] , \mul_b2/fa1_s2_r[15] ,
         \mul_b2/fa1_s2_r[14] , \mul_b2/fa1_s2_r[13] , \mul_b2/fa1_s2_r[12] ,
         \mul_b2/fa1_s1_r[33] , \mul_b2/fa1_s1_r[32] , \mul_b2/fa1_s1_r[31] ,
         \mul_b2/fa1_s1_r[30] , \mul_b2/fa1_s1_r[29] , \mul_b2/fa1_s1_r[28] ,
         \mul_b2/fa1_s1_r[27] , \mul_b2/fa1_s1_r[26] , \mul_b2/fa1_s1_r[25] ,
         \mul_b2/fa1_s1_r[24] , \mul_b2/fa1_s1_r[23] , \mul_b2/fa1_s1_r[22] ,
         \mul_b2/fa1_s1_r[21] , \mul_b2/fa1_s1_r[20] , \mul_b2/fa1_s1_r[19] ,
         \mul_b2/fa1_s1_r[18] , \mul_b2/fa1_s1_r[17] , \mul_b2/fa1_s1_r[16] ,
         \mul_b2/fa1_s1_r[15] , \mul_b2/fa1_s1_r[14] , \mul_b2/fa1_s1_r[13] ,
         \mul_b2/fa1_s1_r[12] , \mul_b2/fa1_s1_r[11] , \mul_b2/fa1_s1_r[10] ,
         \mul_b2/fa1_s1_r[9] , \mul_b2/fa1_s1_r[8] , \mul_b2/fa1_s1_r[7] ,
         \mul_b2/fa1_s1_r[6] , \mul_b2/fa1_s0_r[33] , \mul_b2/fa1_s0_r[32] ,
         \mul_b2/fa1_s0_r[31] , \mul_b2/fa1_s0_r[30] , \mul_b2/fa1_s0_r[29] ,
         \mul_b2/fa1_s0_r[28] , \mul_b2/fa1_s0_r[27] , \mul_b2/fa1_s0_r[26] ,
         \mul_b2/fa1_s0_r[25] , \mul_b2/fa1_s0_r[24] , \mul_b2/fa1_s0_r[23] ,
         \mul_b2/fa1_s0_r[22] , \mul_b2/fa1_s0_r[21] , \mul_b2/fa1_s0_r[20] ,
         \mul_b2/fa1_s0_r[19] , \mul_b2/fa1_s0_r[18] , \mul_b2/fa1_s0_r[17] ,
         \mul_b2/fa1_s0_r[16] , \mul_b2/fa1_s0_r[15] , \mul_b2/fa1_s0_r[14] ,
         \mul_b2/fa1_s0_r[13] , \mul_b2/fa1_s0_r[12] , \mul_b2/fa1_s0_r[11] ,
         \mul_b2/fa1_s0_r[10] , \mul_b2/fa1_s0_r[9] , \mul_b2/fa1_s0_r[8] ,
         \mul_b2/fa1_s0_r[7] , \mul_b2/fa1_s0_r[6] , \mul_b2/fa1_s1[7] ,
         \mul_a1/result_sat[15] , \mul_a1/result_sat[14] ,
         \mul_a1/result_sat[13] , \mul_a1/result_sat[12] ,
         \mul_a1/result_sat[11] , \mul_a1/result_sat[10] ,
         \mul_a1/result_sat[9] , \mul_a1/result_sat[8] ,
         \mul_a1/result_sat[7] , \mul_a1/result_sat[6] ,
         \mul_a1/result_sat[5] , \mul_a1/result_sat[4] ,
         \mul_a1/result_sat[3] , \mul_a1/result_sat[2] ,
         \mul_a1/result_sat[1] , \mul_a1/result_sat[0] , \mul_a1/fa1_c1_r[32] ,
         \mul_a1/fa1_c1_r[31] , \mul_a1/fa1_c1_r[30] , \mul_a1/fa1_c1_r[29] ,
         \mul_a1/fa1_c1_r[28] , \mul_a1/fa1_c1_r[27] , \mul_a1/fa1_c1_r[26] ,
         \mul_a1/fa1_c1_r[25] , \mul_a1/fa1_c1_r[24] , \mul_a1/fa1_c1_r[23] ,
         \mul_a1/fa1_c1_r[22] , \mul_a1/fa1_c1_r[21] , \mul_a1/fa1_c1_r[20] ,
         \mul_a1/fa1_c1_r[19] , \mul_a1/fa1_c1_r[18] , \mul_a1/fa1_c1_r[17] ,
         \mul_a1/fa1_c1_r[16] , \mul_a1/fa1_c1_r[15] , \mul_a1/fa1_c1_r[14] ,
         \mul_a1/fa1_c1_r[13] , \mul_a1/fa1_c1_r[12] , \mul_a1/fa1_c1_r[11] ,
         \mul_a1/fa1_c1_r[10] , \mul_a1/fa1_c1_r[9] , \mul_a1/fa1_c1_r[8] ,
         \mul_a1/fa1_s1_r[33] , \mul_a1/fa1_s1_r[32] , \mul_a1/fa1_s1_r[31] ,
         \mul_a1/fa1_s1_r[30] , \mul_a1/fa1_s1_r[29] , \mul_a1/fa1_s1_r[28] ,
         \mul_a1/fa1_s1_r[27] , \mul_a1/fa1_s1_r[26] , \mul_a1/fa1_s1_r[25] ,
         \mul_a1/fa1_s1_r[24] , \mul_a1/fa1_s1_r[23] , \mul_a1/fa1_s1_r[22] ,
         \mul_a1/fa1_s1_r[21] , \mul_a1/fa1_s1_r[20] , \mul_a1/fa1_s1_r[19] ,
         \mul_a1/fa1_s1_r[18] , \mul_a1/fa1_s1_r[17] , \mul_a1/fa1_s1_r[16] ,
         \mul_a1/fa1_s1_r[15] , \mul_a1/fa1_s1_r[14] , \mul_a1/fa1_s1_r[13] ,
         \mul_a1/fa1_s1_r[12] , \mul_a1/fa1_s1_r[11] , \mul_a1/fa1_s1_r[10] ,
         \mul_a1/fa1_s1_r[9] , \mul_a1/fa1_s1_r[8] , \mul_a1/fa1_s1_r[7] ,
         \mul_a1/fa1_s1_r[6] , \mul_a1/fa1_s0_r[33] , \mul_a1/fa1_s0_r[32] ,
         \mul_a1/fa1_s0_r[31] , \mul_a1/fa1_s0_r[30] , \mul_a1/fa1_s0_r[29] ,
         \mul_a1/fa1_s0_r[28] , \mul_a1/fa1_s0_r[27] , \mul_a1/fa1_s0_r[26] ,
         \mul_a1/fa1_s0_r[25] , \mul_a1/fa1_s0_r[24] , \mul_a1/fa1_s0_r[23] ,
         \mul_a1/fa1_s0_r[22] , \mul_a1/fa1_s0_r[21] , \mul_a1/fa1_s0_r[20] ,
         \mul_a1/fa1_s0_r[19] , \mul_a1/fa1_s0_r[18] , \mul_a1/fa1_s0_r[17] ,
         \mul_a1/fa1_s0_r[16] , \mul_a1/fa1_s0_r[15] , \mul_a1/fa1_s0_r[14] ,
         \mul_a1/fa1_s0_r[13] , \mul_a1/fa1_s0_r[12] , \mul_a1/fa1_s0_r[11] ,
         \mul_a1/fa1_s0_r[10] , \mul_a1/fa1_s0_r[9] , \mul_a1/fa1_s0_r[8] ,
         \mul_a1/fa1_s0_r[7] , \mul_a1/fa1_s0_r[6] , \mul_a1/fa1_c1[23] ,
         \mul_a1/fa1_c1[22] , \mul_a1/fa1_c1[21] , \mul_a1/fa1_c1[20] ,
         \mul_a1/fa1_c1[19] , \mul_a1/fa1_c1[18] , \mul_a1/fa1_c1[17] ,
         \mul_a1/fa1_c1[16] , \mul_a1/fa1_c1[15] , \mul_a1/fa1_c1[14] ,
         \mul_a1/fa1_c1[13] , \mul_a1/fa1_c1[12] , \mul_a1/fa1_c1[11] ,
         \mul_a1/fa1_c1[10] , \mul_a1/fa1_c1[9] , \mul_a1/fa1_c1[8] ,
         \mul_a1/fa1_s1[24] , \mul_a1/fa1_s1[23] , \mul_a1/fa1_s1[22] ,
         \mul_a1/fa1_s1[21] , \mul_a1/fa1_s1[20] , \mul_a1/fa1_s1[19] ,
         \mul_a1/fa1_s1[18] , \mul_a1/fa1_s1[17] , \mul_a1/fa1_s1[16] ,
         \mul_a1/fa1_s1[15] , \mul_a1/fa1_s1[14] , \mul_a1/fa1_s1[13] ,
         \mul_a1/fa1_s1[12] , \mul_a1/fa1_s1[11] , \mul_a1/fa1_s1[10] ,
         \mul_a1/fa1_s1[9] , \mul_a1/fa1_s1[8] , \mul_a2/result_sat[15] ,
         \mul_a2/result_sat[14] , \mul_a2/result_sat[13] ,
         \mul_a2/result_sat[12] , \mul_a2/result_sat[11] ,
         \mul_a2/result_sat[10] , \mul_a2/result_sat[9] ,
         \mul_a2/result_sat[8] , \mul_a2/result_sat[7] ,
         \mul_a2/result_sat[6] , \mul_a2/result_sat[5] ,
         \mul_a2/result_sat[4] , \mul_a2/result_sat[3] ,
         \mul_a2/result_sat[2] , \mul_a2/result_sat[1] ,
         \mul_a2/result_sat[0] , \mul_a2/fa1_s2_r[33] , \mul_a2/fa1_s2_r[32] ,
         \mul_a2/fa1_s2_r[31] , \mul_a2/fa1_s2_r[30] , \mul_a2/fa1_s2_r[29] ,
         \mul_a2/fa1_s2_r[28] , \mul_a2/fa1_s2_r[27] , \mul_a2/fa1_s2_r[26] ,
         \mul_a2/fa1_s2_r[25] , \mul_a2/fa1_s2_r[24] , \mul_a2/fa1_s2_r[23] ,
         \mul_a2/fa1_s2_r[22] , \mul_a2/fa1_s2_r[21] , \mul_a2/fa1_s2_r[20] ,
         \mul_a2/fa1_s2_r[19] , \mul_a2/fa1_s2_r[18] , \mul_a2/fa1_s2_r[17] ,
         \mul_a2/fa1_s2_r[16] , \mul_a2/fa1_s2_r[15] , \mul_a2/fa1_s2_r[14] ,
         \mul_a2/fa1_c1_r[32] , \mul_a2/fa1_c1_r[31] , \mul_a2/fa1_c1_r[30] ,
         \mul_a2/fa1_c1_r[29] , \mul_a2/fa1_c1_r[28] , \mul_a2/fa1_c1_r[27] ,
         \mul_a2/fa1_c1_r[26] , \mul_a2/fa1_c1_r[25] , \mul_a2/fa1_c1_r[24] ,
         \mul_a2/fa1_c1_r[23] , \mul_a2/fa1_c1_r[22] , \mul_a2/fa1_c1_r[21] ,
         \mul_a2/fa1_c1_r[20] , \mul_a2/fa1_c1_r[19] , \mul_a2/fa1_c1_r[18] ,
         \mul_a2/fa1_c1_r[17] , \mul_a2/fa1_c1_r[16] , \mul_a2/fa1_c1_r[15] ,
         \mul_a2/fa1_c1_r[14] , \mul_a2/fa1_c1_r[13] , \mul_a2/fa1_c1_r[12] ,
         \mul_a2/fa1_c1_r[11] , \mul_a2/fa1_c1_r[10] , \mul_a2/fa1_s1_r[25] ,
         \mul_a2/fa1_s1_r[24] , \mul_a2/fa1_s1_r[23] , \mul_a2/fa1_s1_r[22] ,
         \mul_a2/fa1_s1_r[21] , \mul_a2/fa1_s1_r[20] , \mul_a2/fa1_s1_r[19] ,
         \mul_a2/fa1_s1_r[18] , \mul_a2/fa1_s1_r[17] , \mul_a2/fa1_s1_r[16] ,
         \mul_a2/fa1_s1_r[15] , \mul_a2/fa1_s1_r[14] , \mul_a2/fa1_s1_r[13] ,
         \mul_a2/fa1_s1_r[12] , \mul_a2/fa1_s1_r[11] , \mul_a2/fa1_s1_r[10] ,
         \mul_a2/fa1_s1_r[9] , \mul_a2/fa1_c0_r[16] , \mul_a2/fa1_c0_r[15] ,
         \mul_a2/fa1_c0_r[14] , \mul_a2/fa1_c0_r[13] , \mul_a2/fa1_c0_r[12] ,
         \mul_a2/fa1_c0_r[11] , \mul_a2/fa1_c0_r[10] , \mul_a2/fa1_c0_r[9] ,
         \mul_a2/fa1_c0_r[8] , \mul_a2/fa1_c0_r[7] , \mul_a2/fa1_c0_r[6] ,
         \mul_a2/fa1_c0_r[5] , \mul_a2/fa1_c0_r[4] , \mul_a2/fa1_c0_r[3] ,
         \mul_a2/fa1_c0_r[2] , \mul_a2/fa1_s0_r[33] , \mul_a2/fa1_s0_r[32] ,
         \mul_a2/fa1_s0_r[31] , \mul_a2/fa1_s0_r[30] , \mul_a2/fa1_s0_r[29] ,
         \mul_a2/fa1_s0_r[28] , \mul_a2/fa1_s0_r[27] , \mul_a2/fa1_s0_r[26] ,
         \mul_a2/fa1_s0_r[25] , \mul_a2/fa1_s0_r[24] , \mul_a2/fa1_s0_r[23] ,
         \mul_a2/fa1_s0_r[22] , \mul_a2/fa1_s0_r[21] , \mul_a2/fa1_s0_r[20] ,
         \mul_a2/fa1_s0_r[19] , \mul_a2/fa1_s0_r[18] , \mul_a2/fa1_s0_r[17] ,
         \mul_a2/fa1_s0_r[16] , \mul_a2/fa1_s0_r[15] , \mul_a2/fa1_s0_r[14] ,
         \mul_a2/fa1_s0_r[13] , \mul_a2/fa1_s0_r[12] , \mul_a2/fa1_s0_r[11] ,
         \mul_a2/fa1_s0_r[10] , \mul_a2/fa1_s0_r[9] , \mul_a2/fa1_s0_r[8] ,
         \mul_a2/fa1_s0_r[7] , \mul_a2/fa1_s0_r[6] , \mul_a2/fa1_s0_r[5] ,
         \mul_a2/fa1_s0_r[4] , \mul_a2/fa1_s0_r[3] , \mul_a2/fa1_c1[24] ,
         \mul_a2/fa1_c1[23] , \mul_a2/fa1_c1[22] , \mul_a2/fa1_c1[21] ,
         \mul_a2/fa1_c1[20] , \mul_a2/fa1_c1[19] , \mul_a2/fa1_c1[18] ,
         \mul_a2/fa1_c1[17] , \mul_a2/fa1_c1[16] , \mul_a2/fa1_c1[15] ,
         \mul_a2/fa1_c1[14] , \mul_a2/fa1_c1[13] , \mul_a2/fa1_c1[12] ,
         \mul_a2/fa1_c1[11] , \mul_a2/fa1_c1[10] , \mul_a2/fa1_s1[25] ,
         \mul_a2/fa1_s1[24] , \mul_a2/fa1_s1[23] , \mul_a2/fa1_s1[22] ,
         \mul_a2/fa1_s1[21] , \mul_a2/fa1_s1[20] , \mul_a2/fa1_s1[19] ,
         \mul_a2/fa1_s1[18] , \mul_a2/fa1_s1[17] , \mul_a2/fa1_s1[16] ,
         \mul_a2/fa1_s1[15] , \mul_a2/fa1_s1[14] , \mul_a2/fa1_s1[13] ,
         \mul_a2/fa1_s1[12] , \mul_a2/fa1_s1[11] , \mul_a2/fa1_s1[10] ,
         \mul_a2/fa1_c0[16] , \mul_a2/fa1_c0[15] , \mul_a2/fa1_c0[14] ,
         \mul_a2/fa1_c0[13] , \mul_a2/fa1_c0[12] , \mul_a2/fa1_c0[11] ,
         \mul_a2/fa1_c0[10] , \mul_a2/fa1_c0[9] , \mul_a2/fa1_c0[8] ,
         \mul_a2/fa1_c0[7] , \mul_a2/fa1_c0[6] , \mul_a2/fa1_c0[5] ,
         \mul_a2/fa1_c0[4] , \mul_a2/fa1_c0[3] , \mul_a2/fa1_c0[2] ,
         \mul_a2/fa1_s0[28] , \mul_a2/fa1_s0[16] , \mul_a2/fa1_s0[15] ,
         \mul_a2/fa1_s0[14] , \mul_a2/fa1_s0[13] , \mul_a2/fa1_s0[12] ,
         \mul_a2/fa1_s0[11] , \mul_a2/fa1_s0[10] , \mul_a2/fa1_s0[9] ,
         \mul_a2/fa1_s0[8] , \mul_a2/fa1_s0[7] , \mul_a2/fa1_s0[6] ,
         \mul_a2/fa1_s0[5] , \mul_a2/fa1_s0[4] , \mul_a2/fa1_s0[3] ,
         \C50/DATA4_6 , \C50/DATA4_7 , \C50/DATA4_8 , \C50/DATA4_9 ,
         \C50/DATA4_10 , \C50/DATA4_11 , \C50/DATA4_12 , \C50/DATA4_13 ,
         \C50/DATA4_14 , \C50/DATA4_15 , \C50/DATA4_16 , \C50/DATA4_17 ,
         \C50/DATA4_18 , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810;
  wire   [15:0] x_z1;
  wire   [15:0] x_z2;
  wire   [15:0] y_z1;
  wire   [15:0] y_z2;
  wire   [15:0] x_reg2;
  wire   [15:0] p_b0;
  wire   [15:0] p_b1;
  wire   [15:0] p_b2;
  wire   [15:0] p_a1;
  wire   [15:0] p_a2;

  HS65_GS_DFPRQX4 valid_T1_reg ( .D(n1714), .CP(clk), .RN(rst_n), .Q(valid_T1)
         );
  HS65_GS_DFPRQX4 valid_T2_reg ( .D(valid_T1), .CP(clk), .RN(rst_n), .Q(
        valid_T2) );
  HS65_GS_DFPRQX4 valid_T3_reg ( .D(valid_T2), .CP(clk), .RN(rst_n), .Q(
        valid_T3) );
  HS65_GS_DFPRQX4 valid_out_reg ( .D(valid_T3), .CP(clk), .RN(rst_n), .Q(
        valid_out) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[0]  ( .D(\mul_b0/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[0]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[1]  ( .D(\mul_b0/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[1]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[2]  ( .D(\mul_b0/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[2]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[3]  ( .D(\mul_b0/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[3]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[4]  ( .D(\mul_b0/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[4]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[5]  ( .D(\mul_b0/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[5]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[6]  ( .D(\mul_b0/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[6]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[7]  ( .D(\mul_b0/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[7]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[8]  ( .D(\mul_b0/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[8]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[9]  ( .D(\mul_b0/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[9]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[10]  ( .D(\mul_b0/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[10]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[11]  ( .D(\mul_b0/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[11]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[12]  ( .D(\mul_b0/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[12]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[13]  ( .D(\mul_b0/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[13]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[14]  ( .D(\mul_b0/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[14]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[15]  ( .D(\mul_b0/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[15]) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[12]  ( .D(x_z1[0]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[13]  ( .D(x_z1[1]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[14]  ( .D(x_z1[2]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[15]  ( .D(x_z1[3]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[16]  ( .D(x_z1[4]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[17]  ( .D(x_z1[5]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[18]  ( .D(x_z1[6]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[19]  ( .D(x_z1[7]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[20]  ( .D(x_z1[8]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[21]  ( .D(x_z1[9]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[22]  ( .D(x_z1[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[23]  ( .D(x_z1[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[24]  ( .D(x_z1[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[25]  ( .D(x_z1[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[26]  ( .D(x_z1[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[27]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[28]  ( .D(n1713), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[29]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[30]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[31]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[32]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[33]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[8]  ( .D(x_z1[0]), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[9]  ( .D(x_z1[1]), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[10]  ( .D(x_z1[2]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[11]  ( .D(x_z1[3]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[12]  ( .D(x_z1[4]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[13]  ( .D(x_z1[5]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[14]  ( .D(x_z1[6]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[15]  ( .D(x_z1[7]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[16]  ( .D(x_z1[8]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[17]  ( .D(x_z1[9]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[18]  ( .D(x_z1[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[19]  ( .D(x_z1[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[20]  ( .D(x_z1[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[21]  ( .D(x_z1[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[22]  ( .D(x_z1[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[23]  ( .D(n1713), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[24]  ( .D(n1713), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[25]  ( .D(n1713), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[26]  ( .D(n1713), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[27]  ( .D(n1713), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[28]  ( .D(n1713), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[29]  ( .D(n1713), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[30]  ( .D(n1713), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[31]  ( .D(n1713), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[32]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[33]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[5]  ( .D(\mul_b0/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[6]  ( .D(\mul_b0/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[7]  ( .D(\mul_b0/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[8]  ( .D(\mul_b0/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[9]  ( .D(\mul_b0/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[10]  ( .D(\mul_b0/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[11]  ( .D(\mul_b0/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[12]  ( .D(\mul_b0/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[13]  ( .D(\mul_b0/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[14]  ( .D(\mul_b0/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[15]  ( .D(\mul_b0/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[16]  ( .D(\mul_b0/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[17]  ( .D(\mul_b0/fa1_c0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[18]  ( .D(\mul_b0/fa1_c0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[19]  ( .D(\mul_b0/fa1_c0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[20]  ( .D(\mul_b0/fa1_c0[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[6]  ( .D(\mul_b0/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[7]  ( .D(\mul_b0/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[8]  ( .D(\mul_b0/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[9]  ( .D(\mul_b0/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[10]  ( .D(\mul_b0/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[11]  ( .D(\mul_b0/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[12]  ( .D(\mul_b0/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[13]  ( .D(\mul_b0/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[14]  ( .D(\mul_b0/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[15]  ( .D(\mul_b0/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[16]  ( .D(\mul_b0/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[17]  ( .D(\mul_b0/fa1_s0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[18]  ( .D(\mul_b0/fa1_s0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[19]  ( .D(\mul_b0/fa1_s0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[20]  ( .D(\mul_b0/fa1_s0[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[21]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[22]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[23]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[24]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[25]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[26]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[27]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[28]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[29]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[30]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[31]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[32]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[33]  ( .D(\mul_b0/fa1_s0[31] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[0]  ( .D(\mul_b1/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[0]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[1]  ( .D(\mul_b1/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[1]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[2]  ( .D(\mul_b1/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[2]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[3]  ( .D(\mul_b1/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[3]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[4]  ( .D(\mul_b1/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[4]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[5]  ( .D(\mul_b1/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[5]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[6]  ( .D(\mul_b1/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[6]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[7]  ( .D(\mul_b1/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[7]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[8]  ( .D(\mul_b1/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[8]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[9]  ( .D(\mul_b1/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[9]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[10]  ( .D(\mul_b1/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[10]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[11]  ( .D(\mul_b1/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[11]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[12]  ( .D(\mul_b1/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[12]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[13]  ( .D(\mul_b1/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[13]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[14]  ( .D(\mul_b1/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[14]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[15]  ( .D(\mul_b1/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[15]) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[13]  ( .D(\mul_b1/fa1_s0[0] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[14]  ( .D(\mul_b1/fa1_s2[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[15]  ( .D(\mul_b1/fa1_s2[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[16]  ( .D(\mul_b1/fa1_s2[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[17]  ( .D(\mul_b1/fa1_s2[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[18]  ( .D(\mul_b1/fa1_s2[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[19]  ( .D(\mul_b1/fa1_s2[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[20]  ( .D(\mul_b1/fa1_s2[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[21]  ( .D(\mul_b1/fa1_s2[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[22]  ( .D(\mul_b1/fa1_s2[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[23]  ( .D(\mul_b1/fa1_s2[23] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[24]  ( .D(\mul_b1/fa1_s2[24] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[25]  ( .D(\mul_b1/fa1_s2[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[26]  ( .D(\mul_b1/fa1_s2[26] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[27]  ( .D(\mul_b1/fa1_s2[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[28]  ( .D(\mul_b1/fa1_s2[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[29]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[30]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[31]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[32]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[33]  ( .D(\mul_b1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[8]  ( .D(\mul_b1/fa1_c1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[9]  ( .D(\mul_b1/fa1_c1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[10]  ( .D(\mul_b1/fa1_c1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[11]  ( .D(\mul_b1/fa1_c1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[12]  ( .D(\mul_b1/fa1_c1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[13]  ( .D(\mul_b1/fa1_c1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[14]  ( .D(\mul_b1/fa1_c1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[15]  ( .D(\mul_b1/fa1_c1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[16]  ( .D(\mul_b1/fa1_c1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[17]  ( .D(\mul_b1/fa1_c1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[18]  ( .D(\mul_b1/fa1_c1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[19]  ( .D(\mul_b1/fa1_c1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[20]  ( .D(\mul_b1/fa1_c1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[21]  ( .D(\mul_b1/fa1_c1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[22]  ( .D(\mul_b1/fa1_c1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[23]  ( .D(n1712), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[24]  ( .D(n1712), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[25]  ( .D(n1712), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[26]  ( .D(n1712), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[27]  ( .D(n1712), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[28]  ( .D(n1712), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[29]  ( .D(n1712), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[30]  ( .D(n1712), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[31]  ( .D(n1712), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[32]  ( .D(n1712), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[6]  ( .D(\mul_b1/fa1_s0[0] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s1_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[7]  ( .D(\mul_b1/fa1_s0[1] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s1_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[8]  ( .D(\mul_b1/fa1_s1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[9]  ( .D(\mul_b1/fa1_s1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[10]  ( .D(\mul_b1/fa1_s1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[11]  ( .D(\mul_b1/fa1_s1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[12]  ( .D(\mul_b1/fa1_s1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[13]  ( .D(\mul_b1/fa1_s1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[14]  ( .D(\mul_b1/fa1_s1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[15]  ( .D(\mul_b1/fa1_s1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[16]  ( .D(\mul_b1/fa1_s1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[17]  ( .D(\mul_b1/fa1_s1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[18]  ( .D(\mul_b1/fa1_s1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[19]  ( .D(\mul_b1/fa1_s1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[20]  ( .D(\mul_b1/fa1_s1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[21]  ( .D(\mul_b1/fa1_s1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[22]  ( .D(\mul_b1/fa1_s1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[2]  ( .D(n1710), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[2] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[3]  ( .D(n1709), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[3] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[4]  ( .D(\mul_b1/fa1_c0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[5]  ( .D(\mul_b1/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[6]  ( .D(\mul_b1/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[7]  ( .D(\mul_b1/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[8]  ( .D(\mul_b1/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[9]  ( .D(\mul_b1/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[10]  ( .D(\mul_b1/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[11]  ( .D(\mul_b1/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[12]  ( .D(\mul_b1/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[13]  ( .D(\mul_b1/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[14]  ( .D(\mul_b1/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[15]  ( .D(\mul_b1/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[16]  ( .D(\mul_b1/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[17]  ( .D(\mul_b1/fa1_c0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[18]  ( .D(\mul_b1/fa1_c0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[19]  ( .D(n930), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[20]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[21]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[22]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[23]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[24]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[25]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[26]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[27]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[28]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[29]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[30]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[31]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[32]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[3]  ( .D(\mul_b1/fa1_s0[3] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[3] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[4]  ( .D(\mul_b1/fa1_s0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[5]  ( .D(\mul_b1/fa1_s0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[6]  ( .D(\mul_b1/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[7]  ( .D(\mul_b1/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[8]  ( .D(\mul_b1/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[9]  ( .D(\mul_b1/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[10]  ( .D(\mul_b1/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[11]  ( .D(\mul_b1/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[12]  ( .D(\mul_b1/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[13]  ( .D(\mul_b1/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[14]  ( .D(\mul_b1/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[15]  ( .D(\mul_b1/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[16]  ( .D(\mul_b1/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[17]  ( .D(\mul_b1/fa1_s0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[18]  ( .D(\mul_b1/fa1_s0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[19]  ( .D(\mul_b1/fa1_s0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[20]  ( .D(\mul_b1/fa1_s0[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[21]  ( .D(\mul_b1/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[22]  ( .D(\mul_b1/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[23]  ( .D(\mul_b1/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[24]  ( .D(\mul_b1/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[25]  ( .D(\mul_b1/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[26]  ( .D(\mul_b1/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[27]  ( .D(\mul_b1/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[28]  ( .D(\mul_b1/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[29]  ( .D(\mul_b1/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[30]  ( .D(\mul_b1/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[31]  ( .D(\mul_b1/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[32]  ( .D(\mul_b1/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[33]  ( .D(\mul_b1/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[14]  ( .D(\mul_b1/fa1_c2[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[15]  ( .D(\mul_b1/fa1_c2[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[16]  ( .D(\mul_b1/fa1_c2[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[17]  ( .D(\mul_b1/fa1_c2[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[18]  ( .D(\mul_b1/fa1_c2[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[19]  ( .D(\mul_b1/fa1_c2[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[20]  ( .D(\mul_b1/fa1_c2[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[21]  ( .D(\mul_b1/fa1_c2[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[22]  ( .D(\mul_b1/fa1_c2[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[23]  ( .D(\mul_b1/fa1_c2[23] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[24]  ( .D(\mul_b1/fa1_c2[24] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[25]  ( .D(\mul_b1/fa1_c2[25] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[26]  ( .D(\mul_b1/fa1_c2[26] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[27]  ( .D(\mul_b1/fa1_c2[27] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c2_r_reg[28]  ( .D(\mul_b1/fa1_c2[28] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[0]  ( .D(\mul_b2/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[0]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[1]  ( .D(\mul_b2/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[1]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[2]  ( .D(\mul_b2/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[2]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[3]  ( .D(\mul_b2/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[3]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[4]  ( .D(\mul_b2/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[4]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[5]  ( .D(\mul_b2/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[5]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[6]  ( .D(\mul_b2/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[6]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[7]  ( .D(\mul_b2/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[7]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[8]  ( .D(\mul_b2/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[8]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[9]  ( .D(\mul_b2/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[9]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[10]  ( .D(\mul_b2/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[10]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[11]  ( .D(\mul_b2/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[11]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[12]  ( .D(\mul_b2/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[12]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[13]  ( .D(\mul_b2/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[13]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[14]  ( .D(\mul_b2/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[14]) );
  HS65_GS_DFPRQX4 \mul_b2/p_reg[15]  ( .D(\mul_b2/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_b2[15]) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[12]  ( .D(x_reg2[0]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[13]  ( .D(\mul_b2/fa1_s1[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[14]  ( .D(x_reg2[2]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[15]  ( .D(x_reg2[3]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[16]  ( .D(x_reg2[4]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[17]  ( .D(x_reg2[5]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[18]  ( .D(x_reg2[6]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[19]  ( .D(x_reg2[7]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[20]  ( .D(x_reg2[8]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[21]  ( .D(x_reg2[9]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[22]  ( .D(x_reg2[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[23]  ( .D(x_reg2[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[24]  ( .D(x_reg2[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[25]  ( .D(x_reg2[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[26]  ( .D(x_reg2[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[27]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[28]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[29]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[30]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[31]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[32]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s2_r_reg[33]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[6]  ( .D(x_reg2[0]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[7]  ( .D(\mul_b2/fa1_s1[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b2/fa1_s1_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[8]  ( .D(x_reg2[2]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[9]  ( .D(x_reg2[3]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[10]  ( .D(x_reg2[4]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[11]  ( .D(x_reg2[5]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[12]  ( .D(x_reg2[6]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[13]  ( .D(x_reg2[7]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[14]  ( .D(x_reg2[8]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[15]  ( .D(x_reg2[9]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[16]  ( .D(x_reg2[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[17]  ( .D(x_reg2[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[18]  ( .D(x_reg2[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[19]  ( .D(x_reg2[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[20]  ( .D(x_reg2[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[21]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[22]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[23]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[24]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[25]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[26]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[27]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[28]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[29]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[30]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[31]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[32]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s1_r_reg[33]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[6]  ( .D(x_reg2[2]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[7]  ( .D(x_reg2[3]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[8]  ( .D(x_reg2[4]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[9]  ( .D(x_reg2[5]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[10]  ( .D(x_reg2[6]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[11]  ( .D(x_reg2[7]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[12]  ( .D(x_reg2[8]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[13]  ( .D(x_reg2[9]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[14]  ( .D(x_reg2[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[15]  ( .D(x_reg2[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[16]  ( .D(x_reg2[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[17]  ( .D(x_reg2[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[18]  ( .D(x_reg2[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[19]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[20]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[21]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[22]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[23]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[24]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[25]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[26]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[27]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[28]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[29]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[30]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[31]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[32]  ( .D(n1711), .CP(clk), .RN(rst_n), 
        .Q(\mul_b2/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b2/fa1_s0_r_reg[33]  ( .D(x_reg2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b2/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[0]  ( .D(\mul_a1/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[0]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[1]  ( .D(\mul_a1/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[1]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[2]  ( .D(\mul_a1/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[2]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[3]  ( .D(\mul_a1/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[3]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[4]  ( .D(\mul_a1/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[4]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[5]  ( .D(\mul_a1/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[5]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[6]  ( .D(\mul_a1/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[6]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[7]  ( .D(\mul_a1/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[7]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[8]  ( .D(\mul_a1/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[8]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[9]  ( .D(\mul_a1/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[9]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[10]  ( .D(\mul_a1/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[10]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[11]  ( .D(\mul_a1/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[11]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[12]  ( .D(\mul_a1/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[12]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[13]  ( .D(\mul_a1/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[13]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[14]  ( .D(\mul_a1/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[14]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[15]  ( .D(\mul_a1/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[15]) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[8]  ( .D(\mul_a1/fa1_c1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_c1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[9]  ( .D(\mul_a1/fa1_c1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_c1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[10]  ( .D(\mul_a1/fa1_c1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[11]  ( .D(\mul_a1/fa1_c1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[12]  ( .D(\mul_a1/fa1_c1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[13]  ( .D(\mul_a1/fa1_c1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[14]  ( .D(\mul_a1/fa1_c1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[15]  ( .D(\mul_a1/fa1_c1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[16]  ( .D(\mul_a1/fa1_c1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[17]  ( .D(\mul_a1/fa1_c1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[18]  ( .D(\mul_a1/fa1_c1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[19]  ( .D(\mul_a1/fa1_c1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[20]  ( .D(\mul_a1/fa1_c1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[21]  ( .D(\mul_a1/fa1_c1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[22]  ( .D(\mul_a1/fa1_c1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[23]  ( .D(\mul_a1/fa1_c1[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[24]  ( .D(y_z1[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_c1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[25]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_c1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[26]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_c1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[27]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_c1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[28]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_c1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[29]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_c1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[30]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_c1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[31]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_c1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[32]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_c1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[6]  ( .D(y_z1[0]), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[6] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[7]  ( .D(y_z1[1]), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[8]  ( .D(\mul_a1/fa1_s1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[9]  ( .D(\mul_a1/fa1_s1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[10]  ( .D(\mul_a1/fa1_s1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[11]  ( .D(\mul_a1/fa1_s1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[12]  ( .D(\mul_a1/fa1_s1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[13]  ( .D(\mul_a1/fa1_s1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[14]  ( .D(\mul_a1/fa1_s1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[15]  ( .D(\mul_a1/fa1_s1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[16]  ( .D(\mul_a1/fa1_s1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[17]  ( .D(\mul_a1/fa1_s1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[18]  ( .D(\mul_a1/fa1_s1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[19]  ( .D(\mul_a1/fa1_s1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[20]  ( .D(\mul_a1/fa1_s1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[21]  ( .D(\mul_a1/fa1_s1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[22]  ( .D(\mul_a1/fa1_s1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[23]  ( .D(\mul_a1/fa1_s1[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[24]  ( .D(\mul_a1/fa1_s1[24] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[25]  ( .D(n1708), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[26]  ( .D(n1708), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[27]  ( .D(n1708), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[28]  ( .D(n1708), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[29]  ( .D(n1708), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[30]  ( .D(n1708), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[31]  ( .D(n1708), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[32]  ( .D(n1708), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[33]  ( .D(n1708), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[6]  ( .D(\C50/DATA4_6 ), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[7]  ( .D(\C50/DATA4_7 ), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[8]  ( .D(\C50/DATA4_8 ), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[9]  ( .D(\C50/DATA4_9 ), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[10]  ( .D(\C50/DATA4_10 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[11]  ( .D(\C50/DATA4_11 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[12]  ( .D(\C50/DATA4_12 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[13]  ( .D(\C50/DATA4_13 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[14]  ( .D(\C50/DATA4_14 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[15]  ( .D(\C50/DATA4_15 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[16]  ( .D(\C50/DATA4_16 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[17]  ( .D(\C50/DATA4_17 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[18]  ( .D(\C50/DATA4_18 ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[19]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[20]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[21]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[22]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[23]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[24]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[25]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[26]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[27]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[28]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[29]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[30]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[31]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[32]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[33]  ( .D(n1), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[0]  ( .D(\mul_a2/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[0]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[1]  ( .D(\mul_a2/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[1]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[2]  ( .D(\mul_a2/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[2]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[3]  ( .D(\mul_a2/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[3]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[4]  ( .D(\mul_a2/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[4]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[5]  ( .D(\mul_a2/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[5]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[6]  ( .D(\mul_a2/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[6]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[7]  ( .D(\mul_a2/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[7]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[8]  ( .D(\mul_a2/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[8]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[9]  ( .D(\mul_a2/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[9]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[10]  ( .D(\mul_a2/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[10]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[11]  ( .D(\mul_a2/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[11]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[12]  ( .D(\mul_a2/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[12]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[13]  ( .D(\mul_a2/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[13]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[14]  ( .D(\mul_a2/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[14]) );
  HS65_GS_DFPRQX4 \mul_a2/p_reg[15]  ( .D(\mul_a2/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_a2[15]) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[14]  ( .D(y_z2[0]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[15]  ( .D(y_z2[1]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[16]  ( .D(y_z2[2]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[17]  ( .D(y_z2[3]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[18]  ( .D(y_z2[4]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[19]  ( .D(y_z2[5]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[20]  ( .D(y_z2[6]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[21]  ( .D(y_z2[7]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[22]  ( .D(y_z2[8]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[23]  ( .D(y_z2[9]), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[24]  ( .D(y_z2[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[25]  ( .D(y_z2[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[26]  ( .D(y_z2[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[27]  ( .D(y_z2[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[28]  ( .D(y_z2[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[29]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[30]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[31]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[32]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s2_r_reg[33]  ( .D(y_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a2/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[10]  ( .D(\mul_a2/fa1_c1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[11]  ( .D(\mul_a2/fa1_c1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[12]  ( .D(\mul_a2/fa1_c1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[13]  ( .D(\mul_a2/fa1_c1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[14]  ( .D(\mul_a2/fa1_c1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[15]  ( .D(\mul_a2/fa1_c1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[16]  ( .D(\mul_a2/fa1_c1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[17]  ( .D(\mul_a2/fa1_c1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[18]  ( .D(\mul_a2/fa1_c1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[19]  ( .D(\mul_a2/fa1_c1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[20]  ( .D(\mul_a2/fa1_c1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[21]  ( .D(\mul_a2/fa1_c1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[22]  ( .D(\mul_a2/fa1_c1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[23]  ( .D(\mul_a2/fa1_c1[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[24]  ( .D(\mul_a2/fa1_c1[24] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[25]  ( .D(n1707), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[26]  ( .D(n1707), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[27]  ( .D(n1707), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[28]  ( .D(n1707), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[29]  ( .D(n1707), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[30]  ( .D(n1707), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[31]  ( .D(n1707), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c1_r_reg[32]  ( .D(n1707), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_c1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[9]  ( .D(y_z2[0]), .CP(clk), .RN(rst_n), 
        .Q(\mul_a2/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[10]  ( .D(\mul_a2/fa1_s1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[11]  ( .D(\mul_a2/fa1_s1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[12]  ( .D(\mul_a2/fa1_s1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[13]  ( .D(\mul_a2/fa1_s1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[14]  ( .D(\mul_a2/fa1_s1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[15]  ( .D(\mul_a2/fa1_s1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[16]  ( .D(\mul_a2/fa1_s1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[17]  ( .D(\mul_a2/fa1_s1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[18]  ( .D(\mul_a2/fa1_s1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[19]  ( .D(\mul_a2/fa1_s1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[20]  ( .D(\mul_a2/fa1_s1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[21]  ( .D(\mul_a2/fa1_s1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[22]  ( .D(\mul_a2/fa1_s1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[23]  ( .D(\mul_a2/fa1_s1[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[24]  ( .D(\mul_a2/fa1_s1[24] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s1_r_reg[25]  ( .D(\mul_a2/fa1_s1[25] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[2]  ( .D(\mul_a2/fa1_c0[2] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[2] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[3]  ( .D(\mul_a2/fa1_c0[3] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[3] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[4]  ( .D(\mul_a2/fa1_c0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[5]  ( .D(\mul_a2/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[6]  ( .D(\mul_a2/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[7]  ( .D(\mul_a2/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[8]  ( .D(\mul_a2/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[9]  ( .D(\mul_a2/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[10]  ( .D(\mul_a2/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[11]  ( .D(\mul_a2/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[12]  ( .D(\mul_a2/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[13]  ( .D(\mul_a2/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[14]  ( .D(\mul_a2/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[15]  ( .D(\mul_a2/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_c0_r_reg[16]  ( .D(\mul_a2/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[3]  ( .D(\mul_a2/fa1_s0[3] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[3] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[4]  ( .D(\mul_a2/fa1_s0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[5]  ( .D(\mul_a2/fa1_s0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[6]  ( .D(\mul_a2/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[7]  ( .D(\mul_a2/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[8]  ( .D(\mul_a2/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[9]  ( .D(\mul_a2/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a2/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[10]  ( .D(\mul_a2/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[11]  ( .D(\mul_a2/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[12]  ( .D(\mul_a2/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[13]  ( .D(\mul_a2/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[14]  ( .D(\mul_a2/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[15]  ( .D(\mul_a2/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[16]  ( .D(\mul_a2/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[17]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[18]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[19]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[20]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[21]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[22]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[23]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[24]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[25]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[26]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[27]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[28]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[29]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[30]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[31]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[32]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a2/fa1_s0_r_reg[33]  ( .D(\mul_a2/fa1_s0[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a2/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \x_z1_reg[15]  ( .D(n1715), .CP(clk), .RN(rst_n), .Q(
        x_z1[15]) );
  HS65_GS_DFPRQX4 \x_z1_reg[14]  ( .D(n1716), .CP(clk), .RN(rst_n), .Q(
        x_z1[14]) );
  HS65_GS_DFPRQX4 \x_z1_reg[13]  ( .D(n1717), .CP(clk), .RN(rst_n), .Q(
        x_z1[13]) );
  HS65_GS_DFPRQX4 \x_z1_reg[12]  ( .D(n1718), .CP(clk), .RN(rst_n), .Q(
        x_z1[12]) );
  HS65_GS_DFPRQX4 \x_z1_reg[11]  ( .D(n1719), .CP(clk), .RN(rst_n), .Q(
        x_z1[11]) );
  HS65_GS_DFPRQX4 \x_z1_reg[10]  ( .D(n1720), .CP(clk), .RN(rst_n), .Q(
        x_z1[10]) );
  HS65_GS_DFPRQX4 \x_z1_reg[9]  ( .D(n1721), .CP(clk), .RN(rst_n), .Q(x_z1[9])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[8]  ( .D(n1722), .CP(clk), .RN(rst_n), .Q(x_z1[8])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[7]  ( .D(n1723), .CP(clk), .RN(rst_n), .Q(x_z1[7])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[6]  ( .D(n1724), .CP(clk), .RN(rst_n), .Q(x_z1[6])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[5]  ( .D(n1725), .CP(clk), .RN(rst_n), .Q(x_z1[5])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[4]  ( .D(n1726), .CP(clk), .RN(rst_n), .Q(x_z1[4])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[3]  ( .D(n1727), .CP(clk), .RN(rst_n), .Q(x_z1[3])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[2]  ( .D(n1728), .CP(clk), .RN(rst_n), .Q(x_z1[2])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[1]  ( .D(n1729), .CP(clk), .RN(rst_n), .Q(x_z1[1])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[0]  ( .D(n1730), .CP(clk), .RN(rst_n), .Q(x_z1[0])
         );
  HS65_GS_DFPRQX4 \x_z2_reg[15]  ( .D(n1731), .CP(clk), .RN(rst_n), .Q(
        x_z2[15]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[15]  ( .D(n1732), .CP(clk), .RN(rst_n), .Q(
        x_reg2[15]) );
  HS65_GS_DFPRQX4 \x_z2_reg[14]  ( .D(n1733), .CP(clk), .RN(rst_n), .Q(
        x_z2[14]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[14]  ( .D(n1734), .CP(clk), .RN(rst_n), .Q(
        x_reg2[14]) );
  HS65_GS_DFPRQX4 \x_z2_reg[13]  ( .D(n1735), .CP(clk), .RN(rst_n), .Q(
        x_z2[13]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[13]  ( .D(n1736), .CP(clk), .RN(rst_n), .Q(
        x_reg2[13]) );
  HS65_GS_DFPRQX4 \x_z2_reg[12]  ( .D(n1737), .CP(clk), .RN(rst_n), .Q(
        x_z2[12]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[12]  ( .D(n1738), .CP(clk), .RN(rst_n), .Q(
        x_reg2[12]) );
  HS65_GS_DFPRQX4 \x_z2_reg[11]  ( .D(n1739), .CP(clk), .RN(rst_n), .Q(
        x_z2[11]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[11]  ( .D(n1740), .CP(clk), .RN(rst_n), .Q(
        x_reg2[11]) );
  HS65_GS_DFPRQX4 \x_z2_reg[10]  ( .D(n1741), .CP(clk), .RN(rst_n), .Q(
        x_z2[10]) );
  HS65_GS_DFPRQX4 \x_reg2_reg[10]  ( .D(n1742), .CP(clk), .RN(rst_n), .Q(
        x_reg2[10]) );
  HS65_GS_DFPRQX4 \x_z2_reg[9]  ( .D(n1743), .CP(clk), .RN(rst_n), .Q(x_z2[9])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[9]  ( .D(n1744), .CP(clk), .RN(rst_n), .Q(
        x_reg2[9]) );
  HS65_GS_DFPRQX4 \x_z2_reg[8]  ( .D(n1745), .CP(clk), .RN(rst_n), .Q(x_z2[8])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[8]  ( .D(n1746), .CP(clk), .RN(rst_n), .Q(
        x_reg2[8]) );
  HS65_GS_DFPRQX4 \x_z2_reg[7]  ( .D(n1747), .CP(clk), .RN(rst_n), .Q(x_z2[7])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[7]  ( .D(n1748), .CP(clk), .RN(rst_n), .Q(
        x_reg2[7]) );
  HS65_GS_DFPRQX4 \x_z2_reg[6]  ( .D(n1749), .CP(clk), .RN(rst_n), .Q(x_z2[6])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[6]  ( .D(n1750), .CP(clk), .RN(rst_n), .Q(
        x_reg2[6]) );
  HS65_GS_DFPRQX4 \x_z2_reg[5]  ( .D(n1751), .CP(clk), .RN(rst_n), .Q(x_z2[5])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[5]  ( .D(n1752), .CP(clk), .RN(rst_n), .Q(
        x_reg2[5]) );
  HS65_GS_DFPRQX4 \x_z2_reg[4]  ( .D(n1753), .CP(clk), .RN(rst_n), .Q(x_z2[4])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[4]  ( .D(n1754), .CP(clk), .RN(rst_n), .Q(
        x_reg2[4]) );
  HS65_GS_DFPRQX4 \x_z2_reg[3]  ( .D(n1755), .CP(clk), .RN(rst_n), .Q(x_z2[3])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[3]  ( .D(n1756), .CP(clk), .RN(rst_n), .Q(
        x_reg2[3]) );
  HS65_GS_DFPRQX4 \x_z2_reg[2]  ( .D(n1757), .CP(clk), .RN(rst_n), .Q(x_z2[2])
         );
  HS65_GS_DFPRQX4 \x_reg2_reg[2]  ( .D(n1758), .CP(clk), .RN(rst_n), .Q(
        x_reg2[2]) );
  HS65_GS_DFPRQX4 \x_z2_reg[1]  ( .D(n1759), .CP(clk), .RN(rst_n), .Q(
        \mul_b1/fa1_s0[1] ) );
  HS65_GS_DFPRQX4 \x_reg2_reg[1]  ( .D(n1760), .CP(clk), .RN(rst_n), .Q(
        \mul_b2/fa1_s1[7] ) );
  HS65_GS_DFPRQX4 \x_z2_reg[0]  ( .D(n1761), .CP(clk), .RN(rst_n), .Q(
        \mul_b1/fa1_s0[0] ) );
  HS65_GS_DFPRQX4 \x_reg2_reg[0]  ( .D(n1762), .CP(clk), .RN(rst_n), .Q(
        x_reg2[0]) );
  HS65_GS_DFPRQX4 \data_out_reg[15]  ( .D(n1763), .CP(clk), .RN(rst_n), .Q(
        data_out[15]) );
  HS65_GS_DFPRQX4 \y_z1_reg[15]  ( .D(n1764), .CP(clk), .RN(rst_n), .Q(
        y_z1[15]) );
  HS65_GS_DFPRQX4 \y_z2_reg[15]  ( .D(n1765), .CP(clk), .RN(rst_n), .Q(
        y_z2[15]) );
  HS65_GS_DFPRQX4 \data_out_reg[14]  ( .D(n1766), .CP(clk), .RN(rst_n), .Q(
        data_out[14]) );
  HS65_GS_DFPRQX4 \y_z1_reg[14]  ( .D(n1767), .CP(clk), .RN(rst_n), .Q(
        y_z1[14]) );
  HS65_GS_DFPRQX4 \y_z2_reg[14]  ( .D(n1768), .CP(clk), .RN(rst_n), .Q(
        y_z2[14]) );
  HS65_GS_DFPRQX4 \data_out_reg[13]  ( .D(n1769), .CP(clk), .RN(rst_n), .Q(
        data_out[13]) );
  HS65_GS_DFPRQX4 \y_z1_reg[13]  ( .D(n1770), .CP(clk), .RN(rst_n), .Q(
        y_z1[13]) );
  HS65_GS_DFPRQX4 \y_z2_reg[13]  ( .D(n1771), .CP(clk), .RN(rst_n), .Q(
        y_z2[13]) );
  HS65_GS_DFPRQX4 \data_out_reg[12]  ( .D(n1772), .CP(clk), .RN(rst_n), .Q(
        data_out[12]) );
  HS65_GS_DFPRQX4 \y_z1_reg[12]  ( .D(n1773), .CP(clk), .RN(rst_n), .Q(
        y_z1[12]) );
  HS65_GS_DFPRQX4 \y_z2_reg[12]  ( .D(n1774), .CP(clk), .RN(rst_n), .Q(
        y_z2[12]) );
  HS65_GS_DFPRQX4 \data_out_reg[11]  ( .D(n1775), .CP(clk), .RN(rst_n), .Q(
        data_out[11]) );
  HS65_GS_DFPRQX4 \y_z1_reg[11]  ( .D(n1776), .CP(clk), .RN(rst_n), .Q(
        y_z1[11]) );
  HS65_GS_DFPRQX4 \y_z2_reg[11]  ( .D(n1777), .CP(clk), .RN(rst_n), .Q(
        y_z2[11]) );
  HS65_GS_DFPRQX4 \data_out_reg[10]  ( .D(n1778), .CP(clk), .RN(rst_n), .Q(
        data_out[10]) );
  HS65_GS_DFPRQX4 \y_z1_reg[10]  ( .D(n1779), .CP(clk), .RN(rst_n), .Q(
        y_z1[10]) );
  HS65_GS_DFPRQX4 \y_z2_reg[10]  ( .D(n1780), .CP(clk), .RN(rst_n), .Q(
        y_z2[10]) );
  HS65_GS_DFPRQX4 \data_out_reg[9]  ( .D(n1781), .CP(clk), .RN(rst_n), .Q(
        data_out[9]) );
  HS65_GS_DFPRQX4 \y_z1_reg[9]  ( .D(n1782), .CP(clk), .RN(rst_n), .Q(y_z1[9])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[9]  ( .D(n1783), .CP(clk), .RN(rst_n), .Q(y_z2[9])
         );
  HS65_GS_DFPRQX4 \data_out_reg[8]  ( .D(n1784), .CP(clk), .RN(rst_n), .Q(
        data_out[8]) );
  HS65_GS_DFPRQX4 \y_z1_reg[8]  ( .D(n1785), .CP(clk), .RN(rst_n), .Q(y_z1[8])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[8]  ( .D(n1786), .CP(clk), .RN(rst_n), .Q(y_z2[8])
         );
  HS65_GS_DFPRQX4 \data_out_reg[7]  ( .D(n1787), .CP(clk), .RN(rst_n), .Q(
        data_out[7]) );
  HS65_GS_DFPRQX4 \y_z1_reg[7]  ( .D(n1788), .CP(clk), .RN(rst_n), .Q(y_z1[7])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[7]  ( .D(n1789), .CP(clk), .RN(rst_n), .Q(y_z2[7])
         );
  HS65_GS_DFPRQX4 \data_out_reg[6]  ( .D(n1790), .CP(clk), .RN(rst_n), .Q(
        data_out[6]) );
  HS65_GS_DFPRQX4 \y_z1_reg[6]  ( .D(n1791), .CP(clk), .RN(rst_n), .Q(y_z1[6])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[6]  ( .D(n1792), .CP(clk), .RN(rst_n), .Q(y_z2[6])
         );
  HS65_GS_DFPRQX4 \data_out_reg[5]  ( .D(n1793), .CP(clk), .RN(rst_n), .Q(
        data_out[5]) );
  HS65_GS_DFPRQX4 \y_z1_reg[5]  ( .D(n1794), .CP(clk), .RN(rst_n), .Q(y_z1[5])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[5]  ( .D(n1795), .CP(clk), .RN(rst_n), .Q(y_z2[5])
         );
  HS65_GS_DFPRQX4 \data_out_reg[4]  ( .D(n1796), .CP(clk), .RN(rst_n), .Q(
        data_out[4]) );
  HS65_GS_DFPRQX4 \y_z1_reg[4]  ( .D(n1797), .CP(clk), .RN(rst_n), .Q(y_z1[4])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[4]  ( .D(n1798), .CP(clk), .RN(rst_n), .Q(y_z2[4])
         );
  HS65_GS_DFPRQX4 \data_out_reg[3]  ( .D(n1799), .CP(clk), .RN(rst_n), .Q(
        data_out[3]) );
  HS65_GS_DFPRQX4 \y_z1_reg[3]  ( .D(n1800), .CP(clk), .RN(rst_n), .Q(y_z1[3])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[3]  ( .D(n1801), .CP(clk), .RN(rst_n), .Q(y_z2[3])
         );
  HS65_GS_DFPRQX4 \data_out_reg[2]  ( .D(n1802), .CP(clk), .RN(rst_n), .Q(
        data_out[2]) );
  HS65_GS_DFPRQX4 \y_z1_reg[2]  ( .D(n1803), .CP(clk), .RN(rst_n), .Q(y_z1[2])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[2]  ( .D(n1804), .CP(clk), .RN(rst_n), .Q(y_z2[2])
         );
  HS65_GS_DFPRQX4 \data_out_reg[1]  ( .D(n1805), .CP(clk), .RN(rst_n), .Q(
        data_out[1]) );
  HS65_GS_DFPRQX4 \y_z1_reg[1]  ( .D(n1806), .CP(clk), .RN(rst_n), .Q(y_z1[1])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[1]  ( .D(n1807), .CP(clk), .RN(rst_n), .Q(y_z2[1])
         );
  HS65_GS_DFPRQX4 \data_out_reg[0]  ( .D(n1808), .CP(clk), .RN(rst_n), .Q(
        data_out[0]) );
  HS65_GS_DFPRQX4 \y_z1_reg[0]  ( .D(n1809), .CP(clk), .RN(rst_n), .Q(y_z1[0])
         );
  HS65_GS_DFPRQX4 \y_z2_reg[0]  ( .D(n1810), .CP(clk), .RN(rst_n), .Q(y_z2[0])
         );
  HS65_GS_NOR2X3 U3 ( .A(y_z1[15]), .B(n1653), .Z(n1) );
  HS65_GS_NOR2X3 U4 ( .A(n1712), .B(n1348), .Z(n2) );
  HS65_GS_AND2X4 U5 ( .A(\mul_b1/fa1_s0_r[31] ), .B(\mul_b1/fa1_c0_r[30] ), 
        .Z(n5) );
  HS65_GS_NAND2X2 U6 ( .A(\mul_b1/fa1_s0_r[32] ), .B(\mul_b1/fa1_c0_r[31] ), 
        .Z(n199) );
  HS65_GS_OA12X4 U7 ( .A(\mul_b1/fa1_s0_r[32] ), .B(\mul_b1/fa1_c0_r[31] ), 
        .C(n199), .Z(n4) );
  HS65_GSS_XOR2X3 U8 ( .A(\mul_b1/fa1_s2_r[32] ), .B(\mul_b1/fa1_c1_r[31] ), 
        .Z(n3) );
  HS65_GS_FA1X4 U9 ( .A0(n5), .B0(n4), .CI(n3), .CO(n205), .S0(n8) );
  HS65_GSS_XOR2X3 U10 ( .A(\mul_b1/fa1_s2_r[31] ), .B(\mul_b1/fa1_c1_r[30] ), 
        .Z(n193) );
  HS65_GSS_XOR2X3 U11 ( .A(\mul_b1/fa1_s0_r[31] ), .B(\mul_b1/fa1_c0_r[30] ), 
        .Z(n192) );
  HS65_GS_AND2X4 U12 ( .A(\mul_b1/fa1_s0_r[30] ), .B(\mul_b1/fa1_c0_r[29] ), 
        .Z(n191) );
  HS65_GS_AND2X4 U13 ( .A(\mul_b1/fa1_s2_r[31] ), .B(\mul_b1/fa1_c1_r[30] ), 
        .Z(n6) );
  HS65_GS_FA1X4 U14 ( .A0(n8), .B0(n7), .CI(n6), .CO(n202), .S0(n1137) );
  HS65_GS_FA1X4 U15 ( .A0(\mul_b1/fa1_c1_r[28] ), .B0(\mul_b1/fa1_c2_r[28] ), 
        .CI(\mul_b1/fa1_s2_r[29] ), .CO(n187), .S0(n11) );
  HS65_GSS_XOR2X3 U16 ( .A(\mul_b1/fa1_s0_r[29] ), .B(\mul_b1/fa1_c0_r[28] ), 
        .Z(n10) );
  HS65_GS_AND2X4 U17 ( .A(\mul_b1/fa1_s0_r[28] ), .B(\mul_b1/fa1_c0_r[27] ), 
        .Z(n9) );
  HS65_GS_AND2X4 U18 ( .A(\mul_b1/fa1_s0_r[29] ), .B(\mul_b1/fa1_c0_r[28] ), 
        .Z(n190) );
  HS65_GSS_XOR2X3 U19 ( .A(\mul_b1/fa1_s2_r[30] ), .B(\mul_b1/fa1_c1_r[29] ), 
        .Z(n189) );
  HS65_GSS_XOR2X3 U20 ( .A(\mul_b1/fa1_s0_r[30] ), .B(\mul_b1/fa1_c0_r[29] ), 
        .Z(n188) );
  HS65_GS_FA1X4 U21 ( .A0(\mul_b1/fa1_c1_r[27] ), .B0(\mul_b1/fa1_c2_r[27] ), 
        .CI(\mul_b1/fa1_s2_r[28] ), .CO(n184), .S0(n14) );
  HS65_GSS_XOR2X3 U22 ( .A(\mul_b1/fa1_s0_r[28] ), .B(\mul_b1/fa1_c0_r[27] ), 
        .Z(n13) );
  HS65_GS_AND2X4 U23 ( .A(\mul_b1/fa1_s0_r[27] ), .B(\mul_b1/fa1_c0_r[26] ), 
        .Z(n12) );
  HS65_GS_FA1X4 U24 ( .A0(n11), .B0(n10), .CI(n9), .CO(n186), .S0(n182) );
  HS65_GS_FA1X4 U25 ( .A0(\mul_b1/fa1_c1_r[26] ), .B0(\mul_b1/fa1_c2_r[26] ), 
        .CI(\mul_b1/fa1_s2_r[27] ), .CO(n181), .S0(n175) );
  HS65_GSS_XOR2X3 U26 ( .A(\mul_b1/fa1_s0_r[27] ), .B(\mul_b1/fa1_c0_r[26] ), 
        .Z(n174) );
  HS65_GS_AND2X4 U27 ( .A(\mul_b1/fa1_s0_r[26] ), .B(\mul_b1/fa1_c0_r[25] ), 
        .Z(n173) );
  HS65_GS_FA1X4 U28 ( .A0(n14), .B0(n13), .CI(n12), .CO(n183), .S0(n179) );
  HS65_GS_FA1X4 U29 ( .A0(\mul_b1/fa1_c1_r[24] ), .B0(\mul_b1/fa1_c2_r[24] ), 
        .CI(\mul_b1/fa1_s2_r[25] ), .CO(n169), .S0(n163) );
  HS65_GSS_XOR2X3 U30 ( .A(\mul_b1/fa1_s0_r[25] ), .B(\mul_b1/fa1_c0_r[24] ), 
        .Z(n162) );
  HS65_GS_AND2X4 U31 ( .A(\mul_b1/fa1_s0_r[24] ), .B(\mul_b1/fa1_c0_r[23] ), 
        .Z(n161) );
  HS65_GS_AND2X4 U32 ( .A(\mul_b1/fa1_s0_r[25] ), .B(\mul_b1/fa1_c0_r[24] ), 
        .Z(n172) );
  HS65_GSS_XOR2X3 U33 ( .A(\mul_b1/fa1_s0_r[26] ), .B(\mul_b1/fa1_c0_r[25] ), 
        .Z(n170) );
  HS65_GS_FA1X4 U34 ( .A0(\mul_b1/fa1_c1_r[22] ), .B0(\mul_b1/fa1_c2_r[22] ), 
        .CI(\mul_b1/fa1_s2_r[23] ), .CO(n157), .S0(n151) );
  HS65_GSS_XOR2X3 U35 ( .A(\mul_b1/fa1_s0_r[23] ), .B(\mul_b1/fa1_c0_r[22] ), 
        .Z(n150) );
  HS65_GS_AND2X4 U36 ( .A(\mul_b1/fa1_s0_r[23] ), .B(\mul_b1/fa1_c0_r[22] ), 
        .Z(n160) );
  HS65_GSS_XOR2X3 U37 ( .A(\mul_b1/fa1_s0_r[24] ), .B(\mul_b1/fa1_c0_r[23] ), 
        .Z(n158) );
  HS65_GS_FA1X4 U38 ( .A0(\mul_b1/fa1_c1_r[20] ), .B0(\mul_b1/fa1_c2_r[20] ), 
        .CI(\mul_b1/fa1_s2_r[21] ), .CO(n145), .S0(n17) );
  HS65_GS_FA1X4 U39 ( .A0(\mul_b1/fa1_s0_r[21] ), .B0(\mul_b1/fa1_s1_r[21] ), 
        .CI(\mul_b1/fa1_c0_r[20] ), .CO(n147), .S0(n15) );
  HS65_GS_FA1X4 U40 ( .A0(\mul_b1/fa1_s0_r[22] ), .B0(\mul_b1/fa1_s1_r[22] ), 
        .CI(\mul_b1/fa1_c0_r[21] ), .CO(n149), .S0(n146) );
  HS65_GS_FA1X4 U41 ( .A0(\mul_b1/fa1_c1_r[19] ), .B0(\mul_b1/fa1_c2_r[19] ), 
        .CI(\mul_b1/fa1_s2_r[20] ), .CO(n140), .S0(n134) );
  HS65_GS_FA1X4 U42 ( .A0(\mul_b1/fa1_s0_r[20] ), .B0(\mul_b1/fa1_s1_r[20] ), 
        .CI(\mul_b1/fa1_c0_r[19] ), .CO(n16), .S0(n132) );
  HS65_GS_FA1X4 U43 ( .A0(n17), .B0(n16), .CI(n15), .CO(n144), .S0(n138) );
  HS65_GS_FA1X4 U44 ( .A0(\mul_b1/fa1_c1_r[16] ), .B0(\mul_b1/fa1_c2_r[16] ), 
        .CI(\mul_b1/fa1_s2_r[17] ), .CO(n122), .S0(n116) );
  HS65_GS_FA1X4 U45 ( .A0(\mul_b1/fa1_s0_r[17] ), .B0(\mul_b1/fa1_s1_r[17] ), 
        .CI(\mul_b1/fa1_c0_r[16] ), .CO(n124), .S0(n114) );
  HS65_GS_AND2X4 U46 ( .A(\mul_b1/fa1_c1_r[13] ), .B(\mul_b1/fa1_s2_r[14] ), 
        .Z(n20) );
  HS65_GSS_XOR2X3 U47 ( .A(\mul_b1/fa1_c1_r[13] ), .B(\mul_b1/fa1_s2_r[14] ), 
        .Z(n98) );
  HS65_GS_FA1X4 U48 ( .A0(\mul_b1/fa1_s0_r[14] ), .B0(\mul_b1/fa1_s1_r[14] ), 
        .CI(\mul_b1/fa1_c0_r[13] ), .CO(n105), .S0(n97) );
  HS65_GS_FA1X4 U49 ( .A0(n20), .B0(n19), .CI(n18), .CO(n1562), .S0(n1558) );
  HS65_GS_FA1X4 U50 ( .A0(\mul_b1/fa1_s0_r[13] ), .B0(\mul_b1/fa1_s1_r[13] ), 
        .CI(\mul_b1/fa1_c0_r[12] ), .CO(n96), .S0(n100) );
  HS65_GSS_XOR2X3 U51 ( .A(\mul_b1/fa1_s2_r[13] ), .B(\mul_b1/fa1_c1_r[12] ), 
        .Z(n99) );
  HS65_GS_PAOI2X1 U52 ( .A(\mul_b1/fa1_s1_r[11] ), .B(\mul_b1/fa1_c0_r[10] ), 
        .P(\mul_b1/fa1_s0_r[11] ), .Z(n21) );
  HS65_GS_IVX2 U53 ( .A(\mul_b1/fa1_c1_r[11] ), .Z(n22) );
  HS65_GS_MUXI21X2 U54 ( .D0(\mul_b1/fa1_c1_r[11] ), .D1(n22), .S0(n21), .Z(
        n80) );
  HS65_GS_FA1X4 U55 ( .A0(\mul_b1/fa1_s0_r[12] ), .B0(\mul_b1/fa1_s1_r[12] ), 
        .CI(\mul_b1/fa1_c0_r[11] ), .CO(n101), .S0(n79) );
  HS65_GS_NAND2X2 U56 ( .A(n80), .B(n79), .Z(n78) );
  HS65_GS_NAND2X2 U57 ( .A(n21), .B(n78), .Z(n24) );
  HS65_GS_NAND2X2 U58 ( .A(n22), .B(n78), .Z(n23) );
  HS65_GS_NAND2X2 U59 ( .A(n24), .B(n23), .Z(n95) );
  HS65_GSS_XOR2X3 U60 ( .A(n93), .B(n95), .Z(n92) );
  HS65_GSS_XOR3X2 U61 ( .A(\mul_b1/fa1_s1_r[10] ), .B(\mul_b1/fa1_c0_r[9] ), 
        .C(\mul_b1/fa1_s0_r[10] ), .Z(n34) );
  HS65_GS_PAO2X4 U62 ( .A(\mul_b1/fa1_s0_r[9] ), .B(\mul_b1/fa1_c0_r[8] ), .P(
        \mul_b1/fa1_s1_r[9] ), .Z(n25) );
  HS65_GSS_XOR2X3 U63 ( .A(\mul_b1/fa1_c1_r[9] ), .B(n25), .Z(n35) );
  HS65_GS_NAND2X2 U64 ( .A(n34), .B(n35), .Z(n33) );
  HS65_GS_NAND2X2 U65 ( .A(\mul_b1/fa1_c1_r[9] ), .B(n25), .Z(n26) );
  HS65_GS_NAND2X2 U66 ( .A(n33), .B(n26), .Z(n31) );
  HS65_GS_IVX2 U67 ( .A(n31), .Z(n29) );
  HS65_GS_PAOI2X1 U68 ( .A(\mul_b1/fa1_s1_r[10] ), .B(\mul_b1/fa1_c0_r[9] ), 
        .P(\mul_b1/fa1_s0_r[10] ), .Z(n75) );
  HS65_GSS_XNOR2X3 U69 ( .A(\mul_b1/fa1_c1_r[10] ), .B(n75), .Z(n28) );
  HS65_GSS_XOR3X2 U70 ( .A(\mul_b1/fa1_s1_r[11] ), .B(\mul_b1/fa1_c0_r[10] ), 
        .C(\mul_b1/fa1_s0_r[11] ), .Z(n27) );
  HS65_GS_NAND2X2 U71 ( .A(n27), .B(n28), .Z(n85) );
  HS65_GS_OAI21X2 U72 ( .A(n28), .B(n27), .C(n85), .Z(n30) );
  HS65_GS_NOR2X2 U73 ( .A(n29), .B(n30), .Z(n84) );
  HS65_GSS_XOR2X3 U74 ( .A(n31), .B(n30), .Z(n74) );
  HS65_GS_IVX2 U75 ( .A(\mul_b1/fa1_c1_r[8] ), .Z(n32) );
  HS65_GS_PAOI2X1 U76 ( .A(\mul_b1/fa1_c0_r[7] ), .B(\mul_b1/fa1_s1_r[8] ), 
        .P(\mul_b1/fa1_s0_r[8] ), .Z(n59) );
  HS65_GS_NOR2X2 U77 ( .A(n32), .B(n59), .Z(n70) );
  HS65_GS_OAI21X2 U78 ( .A(n35), .B(n34), .C(n33), .Z(n68) );
  HS65_GSS_XNOR2X3 U79 ( .A(n70), .B(n68), .Z(n66) );
  HS65_GSS_XNOR3X2 U80 ( .A(\mul_b1/fa1_c0_r[7] ), .B(\mul_b1/fa1_s1_r[8] ), 
        .C(\mul_b1/fa1_s0_r[8] ), .Z(n38) );
  HS65_GS_IVX2 U81 ( .A(n38), .Z(n37) );
  HS65_GS_PAOI2X1 U82 ( .A(\mul_b1/fa1_s1_r[7] ), .B(\mul_b1/fa1_c0_r[6] ), 
        .P(\mul_b1/fa1_s0_r[7] ), .Z(n39) );
  HS65_GS_IVX2 U83 ( .A(n39), .Z(n36) );
  HS65_GS_NAND2X2 U84 ( .A(n37), .B(n36), .Z(n64) );
  HS65_GSS_XNOR3X2 U85 ( .A(\mul_b1/fa1_s1_r[7] ), .B(\mul_b1/fa1_c0_r[6] ), 
        .C(\mul_b1/fa1_s0_r[7] ), .Z(n51) );
  HS65_GS_PAOI2X1 U86 ( .A(\mul_b1/fa1_c0_r[5] ), .B(\mul_b1/fa1_s1_r[6] ), 
        .P(\mul_b1/fa1_s0_r[6] ), .Z(n52) );
  HS65_GS_NOR2X2 U87 ( .A(n51), .B(n52), .Z(n58) );
  HS65_GSS_XOR2X3 U88 ( .A(n39), .B(n38), .Z(n57) );
  HS65_GSS_XNOR3X2 U89 ( .A(\mul_b1/fa1_c0_r[5] ), .B(\mul_b1/fa1_s1_r[6] ), 
        .C(\mul_b1/fa1_s0_r[6] ), .Z(n50) );
  HS65_GS_IVX2 U90 ( .A(n50), .Z(n48) );
  HS65_GS_NAND2X2 U91 ( .A(\mul_b1/fa1_c0_r[3] ), .B(\mul_b1/fa1_s0_r[4] ), 
        .Z(n40) );
  HS65_GSS_XNOR2X3 U92 ( .A(\mul_b1/fa1_c0_r[4] ), .B(\mul_b1/fa1_s0_r[5] ), 
        .Z(n41) );
  HS65_GS_NOR2X2 U93 ( .A(n40), .B(n41), .Z(n47) );
  HS65_GS_IVX2 U94 ( .A(n41), .Z(n45) );
  HS65_GSS_XNOR2X3 U95 ( .A(\mul_b1/fa1_c0_r[3] ), .B(\mul_b1/fa1_s0_r[4] ), 
        .Z(n43) );
  HS65_GS_NAND2X2 U96 ( .A(\mul_b1/fa1_c0_r[2] ), .B(\mul_b1/fa1_s0_r[3] ), 
        .Z(n42) );
  HS65_GS_NOR2X2 U97 ( .A(n43), .B(n42), .Z(n44) );
  HS65_GS_AND2X4 U98 ( .A(n45), .B(n44), .Z(n46) );
  HS65_GS_PAO2X4 U99 ( .A(n48), .B(n47), .P(n46), .Z(n55) );
  HS65_GS_NAND2X2 U100 ( .A(\mul_b1/fa1_c0_r[4] ), .B(\mul_b1/fa1_s0_r[5] ), 
        .Z(n49) );
  HS65_GS_NOR2X2 U101 ( .A(n50), .B(n49), .Z(n54) );
  HS65_GSS_XOR2X3 U102 ( .A(n52), .B(n51), .Z(n53) );
  HS65_GS_PAO2X4 U103 ( .A(n55), .B(n54), .P(n53), .Z(n56) );
  HS65_GS_PAOI2X1 U104 ( .A(n58), .B(n57), .P(n56), .Z(n63) );
  HS65_GSS_XNOR2X3 U105 ( .A(\mul_b1/fa1_c1_r[8] ), .B(n59), .Z(n61) );
  HS65_GSS_XOR3X2 U106 ( .A(\mul_b1/fa1_s0_r[9] ), .B(\mul_b1/fa1_c0_r[8] ), 
        .C(\mul_b1/fa1_s1_r[9] ), .Z(n60) );
  HS65_GS_NAND2X2 U107 ( .A(n60), .B(n61), .Z(n67) );
  HS65_GS_OAI21X2 U108 ( .A(n61), .B(n60), .C(n67), .Z(n62) );
  HS65_GS_PAOI2X1 U109 ( .A(n64), .B(n63), .P(n62), .Z(n65) );
  HS65_GS_NAND2X2 U110 ( .A(n66), .B(n65), .Z(n73) );
  HS65_GS_IVX2 U111 ( .A(n67), .Z(n71) );
  HS65_GS_IVX2 U112 ( .A(n68), .Z(n69) );
  HS65_GS_OAI21X2 U113 ( .A(n71), .B(n70), .C(n69), .Z(n72) );
  HS65_GS_PAOI2X1 U114 ( .A(n74), .B(n73), .P(n72), .Z(n83) );
  HS65_GS_IVX2 U115 ( .A(\mul_b1/fa1_c1_r[10] ), .Z(n76) );
  HS65_GS_NOR2X2 U116 ( .A(n76), .B(n75), .Z(n88) );
  HS65_GS_IVX2 U117 ( .A(n88), .Z(n77) );
  HS65_GS_NAND2X2 U118 ( .A(n77), .B(n85), .Z(n81) );
  HS65_GS_OAI21X2 U119 ( .A(n80), .B(n79), .C(n78), .Z(n86) );
  HS65_GSS_XNOR2X3 U120 ( .A(n81), .B(n86), .Z(n82) );
  HS65_GS_PAOI2X1 U121 ( .A(n84), .B(n83), .P(n82), .Z(n91) );
  HS65_GS_IVX2 U122 ( .A(n85), .Z(n89) );
  HS65_GS_IVX2 U123 ( .A(n86), .Z(n87) );
  HS65_GS_OAI21X2 U124 ( .A(n89), .B(n88), .C(n87), .Z(n90) );
  HS65_GS_PAOI2X1 U125 ( .A(n92), .B(n91), .P(n90), .Z(n1124) );
  HS65_GS_IVX2 U126 ( .A(n93), .Z(n94) );
  HS65_GS_NOR2X2 U127 ( .A(n95), .B(n94), .Z(n1123) );
  HS65_GS_AND2X4 U128 ( .A(\mul_b1/fa1_s2_r[13] ), .B(\mul_b1/fa1_c1_r[12] ), 
        .Z(n104) );
  HS65_GS_FA1X4 U129 ( .A0(n98), .B0(n97), .CI(n96), .CO(n18), .S0(n103) );
  HS65_GS_FA1X4 U130 ( .A0(n101), .B0(n100), .CI(n99), .CO(n102), .S0(n93) );
  HS65_GS_PAO2X4 U131 ( .A(n1124), .B(n1123), .P(n1146), .Z(n1557) );
  HS65_GS_FA1X4 U132 ( .A0(n104), .B0(n103), .CI(n102), .CO(n1556), .S0(n1146)
         );
  HS65_GS_FA1X4 U133 ( .A0(\mul_b1/fa1_c1_r[14] ), .B0(\mul_b1/fa1_c2_r[14] ), 
        .CI(\mul_b1/fa1_s2_r[15] ), .CO(n110), .S0(n106) );
  HS65_GS_FA1X4 U134 ( .A0(n107), .B0(n106), .CI(n105), .CO(n109), .S0(n19) );
  HS65_GS_FA1X4 U135 ( .A0(\mul_b1/fa1_s0_r[15] ), .B0(\mul_b1/fa1_s1_r[15] ), 
        .CI(\mul_b1/fa1_c0_r[14] ), .CO(n112), .S0(n107) );
  HS65_GS_FA1X4 U136 ( .A0(\mul_b1/fa1_s0_r[16] ), .B0(\mul_b1/fa1_s1_r[16] ), 
        .CI(\mul_b1/fa1_c0_r[15] ), .CO(n115), .S0(n111) );
  HS65_GS_FA1X4 U137 ( .A0(n110), .B0(n109), .CI(n108), .CO(n1565), .S0(n1560)
         );
  HS65_GS_FA1X4 U138 ( .A0(\mul_b1/fa1_c1_r[15] ), .B0(\mul_b1/fa1_c2_r[15] ), 
        .CI(\mul_b1/fa1_s2_r[16] ), .CO(n119), .S0(n113) );
  HS65_GS_FA1X4 U139 ( .A0(n113), .B0(n112), .CI(n111), .CO(n118), .S0(n108)
         );
  HS65_GS_FA1X4 U140 ( .A0(n116), .B0(n115), .CI(n114), .CO(n121), .S0(n117)
         );
  HS65_GS_FA1X4 U141 ( .A0(n119), .B0(n118), .CI(n117), .CO(n1569), .S0(n1564)
         );
  HS65_GS_FA1X4 U142 ( .A0(n122), .B0(n121), .CI(n120), .CO(n1574), .S0(n1568)
         );
  HS65_GS_FA1X4 U143 ( .A0(\mul_b1/fa1_c1_r[17] ), .B0(\mul_b1/fa1_c2_r[17] ), 
        .CI(\mul_b1/fa1_s2_r[18] ), .CO(n128), .S0(n125) );
  HS65_GS_FA1X4 U144 ( .A0(n125), .B0(n124), .CI(n123), .CO(n127), .S0(n120)
         );
  HS65_GS_FA1X4 U145 ( .A0(\mul_b1/fa1_s0_r[18] ), .B0(\mul_b1/fa1_s1_r[18] ), 
        .CI(\mul_b1/fa1_c0_r[17] ), .CO(n130), .S0(n123) );
  HS65_GS_FA1X4 U146 ( .A0(\mul_b1/fa1_s0_r[19] ), .B0(\mul_b1/fa1_s1_r[19] ), 
        .CI(\mul_b1/fa1_c0_r[18] ), .CO(n133), .S0(n129) );
  HS65_GS_FA1X4 U147 ( .A0(n128), .B0(n127), .CI(n126), .CO(n1577), .S0(n1572)
         );
  HS65_GS_FA1X4 U148 ( .A0(\mul_b1/fa1_c1_r[18] ), .B0(\mul_b1/fa1_c2_r[18] ), 
        .CI(\mul_b1/fa1_s2_r[19] ), .CO(n137), .S0(n131) );
  HS65_GS_FA1X4 U149 ( .A0(n131), .B0(n130), .CI(n129), .CO(n136), .S0(n126)
         );
  HS65_GS_FA1X4 U150 ( .A0(n134), .B0(n133), .CI(n132), .CO(n139), .S0(n135)
         );
  HS65_GS_FA1X4 U151 ( .A0(n137), .B0(n136), .CI(n135), .CO(n1149), .S0(n1576)
         );
  HS65_GS_NAND2X2 U152 ( .A(n1148), .B(n1149), .Z(n142) );
  HS65_GS_FA1X4 U153 ( .A0(n140), .B0(n139), .CI(n138), .CO(n1582), .S0(n1153)
         );
  HS65_GS_IVX2 U154 ( .A(n1153), .Z(n141) );
  HS65_GS_NOR2X2 U155 ( .A(n1148), .B(n1149), .Z(n1147) );
  HS65_GS_AOI12X2 U156 ( .A(n142), .B(n141), .C(n1147), .Z(n1581) );
  HS65_GS_FA1X4 U157 ( .A0(n145), .B0(n144), .CI(n143), .CO(n1586), .S0(n1580)
         );
  HS65_GS_FA1X4 U158 ( .A0(\mul_b1/fa1_c1_r[21] ), .B0(\mul_b1/fa1_c2_r[21] ), 
        .CI(\mul_b1/fa1_s2_r[22] ), .CO(n154), .S0(n148) );
  HS65_GS_FA1X4 U159 ( .A0(n148), .B0(n147), .CI(n146), .CO(n153), .S0(n143)
         );
  HS65_GS_FA1X4 U160 ( .A0(n151), .B0(n150), .CI(n149), .CO(n156), .S0(n152)
         );
  HS65_GS_FA1X4 U161 ( .A0(n154), .B0(n153), .CI(n152), .CO(n1589), .S0(n1584)
         );
  HS65_GS_FA1X4 U162 ( .A0(n157), .B0(n156), .CI(n155), .CO(n1594), .S0(n1588)
         );
  HS65_GS_FA1X4 U163 ( .A0(\mul_b1/fa1_c1_r[23] ), .B0(\mul_b1/fa1_c2_r[23] ), 
        .CI(\mul_b1/fa1_s2_r[24] ), .CO(n166), .S0(n159) );
  HS65_GS_FA1X4 U164 ( .A0(n160), .B0(n159), .CI(n158), .CO(n165), .S0(n155)
         );
  HS65_GS_FA1X4 U165 ( .A0(n163), .B0(n162), .CI(n161), .CO(n168), .S0(n164)
         );
  HS65_GS_FA1X4 U166 ( .A0(n166), .B0(n165), .CI(n164), .CO(n1597), .S0(n1592)
         );
  HS65_GS_FA1X4 U167 ( .A0(n169), .B0(n168), .CI(n167), .CO(n1602), .S0(n1596)
         );
  HS65_GS_FA1X4 U168 ( .A0(\mul_b1/fa1_c1_r[25] ), .B0(\mul_b1/fa1_c2_r[25] ), 
        .CI(\mul_b1/fa1_s2_r[26] ), .CO(n178), .S0(n171) );
  HS65_GS_FA1X4 U169 ( .A0(n172), .B0(n171), .CI(n170), .CO(n177), .S0(n167)
         );
  HS65_GS_FA1X4 U170 ( .A0(n175), .B0(n174), .CI(n173), .CO(n180), .S0(n176)
         );
  HS65_GS_FA1X4 U171 ( .A0(n178), .B0(n177), .CI(n176), .CO(n1605), .S0(n1600)
         );
  HS65_GS_FA1X4 U172 ( .A0(n181), .B0(n180), .CI(n179), .CO(n1134), .S0(n1604)
         );
  HS65_GS_FA1X4 U173 ( .A0(n184), .B0(n183), .CI(n182), .CO(n1127), .S0(n1132)
         );
  HS65_GS_FA1X4 U174 ( .A0(n187), .B0(n186), .CI(n185), .CO(n1131), .S0(n1125)
         );
  HS65_GS_AND2X4 U175 ( .A(\mul_b1/fa1_c1_r[29] ), .B(\mul_b1/fa1_s2_r[30] ), 
        .Z(n196) );
  HS65_GS_FA1X4 U176 ( .A0(n190), .B0(n189), .CI(n188), .CO(n195), .S0(n185)
         );
  HS65_GS_FA1X4 U177 ( .A0(n193), .B0(n192), .CI(n191), .CO(n7), .S0(n194) );
  HS65_GS_FA1X4 U178 ( .A0(n196), .B0(n195), .CI(n194), .CO(n1135), .S0(n1129)
         );
  HS65_GS_AND2X4 U179 ( .A(\mul_b1/fa1_c1_r[31] ), .B(\mul_b1/fa1_s2_r[32] ), 
        .Z(n197) );
  HS65_GSS_XOR3X2 U180 ( .A(n198), .B(\mul_b1/fa1_c0_r[32] ), .C(n197), .Z(
        n201) );
  HS65_GS_IVX2 U181 ( .A(n199), .Z(n200) );
  HS65_GSS_XOR3X2 U182 ( .A(n202), .B(n201), .C(n200), .Z(n203) );
  HS65_GSS_XOR3X2 U183 ( .A(\mul_b1/fa1_s0_r[33] ), .B(\mul_b1/fa1_c1_r[32] ), 
        .C(n203), .Z(n204) );
  HS65_GSS_XOR3X2 U184 ( .A(n205), .B(\mul_b1/fa1_s2_r[33] ), .C(n204), .Z(
        \mul_b1/result_sat[15] ) );
  HS65_GS_NAND2X2 U185 ( .A(\mul_a2/fa1_c1_r[31] ), .B(\mul_a2/fa1_s2_r[32] ), 
        .Z(n419) );
  HS65_GS_OA12X4 U186 ( .A(\mul_a2/fa1_c1_r[31] ), .B(\mul_a2/fa1_s2_r[32] ), 
        .C(n419), .Z(n206) );
  HS65_GS_AND2X4 U187 ( .A(n206), .B(\mul_a2/fa1_s0_r[32] ), .Z(n418) );
  HS65_GS_AND2X4 U188 ( .A(\mul_a2/fa1_c1_r[30] ), .B(\mul_a2/fa1_s2_r[31] ), 
        .Z(n209) );
  HS65_GSS_XOR2X3 U189 ( .A(\mul_a2/fa1_s0_r[32] ), .B(n206), .Z(n208) );
  HS65_GSS_XOR2X3 U190 ( .A(\mul_a2/fa1_c1_r[30] ), .B(\mul_a2/fa1_s2_r[31] ), 
        .Z(n408) );
  HS65_GS_AND2X4 U191 ( .A(n408), .B(\mul_a2/fa1_s0_r[31] ), .Z(n207) );
  HS65_GS_FA1X4 U192 ( .A0(n209), .B0(n208), .CI(n207), .CO(n416), .S0(n210)
         );
  HS65_GS_IVX2 U193 ( .A(n210), .Z(n883) );
  HS65_GSS_XOR2X3 U194 ( .A(\mul_a2/fa1_s2_r[29] ), .B(\mul_a2/fa1_c1_r[28] ), 
        .Z(n403) );
  HS65_GS_NAND2X2 U195 ( .A(n403), .B(\mul_a2/fa1_s0_r[29] ), .Z(n213) );
  HS65_GS_IVX2 U196 ( .A(n213), .Z(n211) );
  HS65_GS_AND2X4 U197 ( .A(\mul_a2/fa1_s2_r[29] ), .B(\mul_a2/fa1_c1_r[28] ), 
        .Z(n402) );
  HS65_GSS_XOR2X3 U198 ( .A(\mul_a2/fa1_c1_r[29] ), .B(\mul_a2/fa1_s2_r[30] ), 
        .Z(n409) );
  HS65_GSS_XOR2X3 U199 ( .A(n409), .B(\mul_a2/fa1_s0_r[30] ), .Z(n407) );
  HS65_GS_IVX2 U200 ( .A(n407), .Z(n406) );
  HS65_GS_OAI21X2 U201 ( .A(n211), .B(n402), .C(n407), .Z(n886) );
  HS65_GSS_XOR2X3 U202 ( .A(\mul_a2/fa1_s2_r[28] ), .B(\mul_a2/fa1_c1_r[27] ), 
        .Z(n218) );
  HS65_GS_NAND2X2 U203 ( .A(n218), .B(\mul_a2/fa1_s0_r[28] ), .Z(n217) );
  HS65_GS_IVX2 U204 ( .A(n217), .Z(n215) );
  HS65_GS_AND2X4 U205 ( .A(\mul_a2/fa1_s2_r[28] ), .B(\mul_a2/fa1_c1_r[27] ), 
        .Z(n214) );
  HS65_GS_AOI12X2 U206 ( .A(\mul_a2/fa1_s0_r[28] ), .B(n218), .C(n214), .Z(
        n212) );
  HS65_GS_IVX2 U207 ( .A(n212), .Z(n401) );
  HS65_GS_OAI21X2 U208 ( .A(n403), .B(\mul_a2/fa1_s0_r[29] ), .C(n213), .Z(
        n400) );
  HS65_GS_NAND2X2 U209 ( .A(n401), .B(n400), .Z(n399) );
  HS65_GS_OAI21X2 U210 ( .A(n215), .B(n214), .C(n399), .Z(n877) );
  HS65_GSS_XOR2X3 U211 ( .A(\mul_a2/fa1_s2_r[27] ), .B(\mul_a2/fa1_c1_r[26] ), 
        .Z(n390) );
  HS65_GS_NAND2X2 U212 ( .A(n390), .B(\mul_a2/fa1_s0_r[27] ), .Z(n389) );
  HS65_GS_IVX2 U213 ( .A(n389), .Z(n220) );
  HS65_GS_AND2X4 U214 ( .A(\mul_a2/fa1_s2_r[27] ), .B(\mul_a2/fa1_c1_r[26] ), 
        .Z(n219) );
  HS65_GS_AOI12X2 U215 ( .A(\mul_a2/fa1_s0_r[27] ), .B(n390), .C(n219), .Z(
        n216) );
  HS65_GS_IVX2 U216 ( .A(n216), .Z(n398) );
  HS65_GS_OAI21X2 U217 ( .A(n218), .B(\mul_a2/fa1_s0_r[28] ), .C(n217), .Z(
        n397) );
  HS65_GS_NAND2X2 U218 ( .A(n398), .B(n397), .Z(n396) );
  HS65_GS_OAI21X2 U219 ( .A(n220), .B(n219), .C(n396), .Z(n880) );
  HS65_GS_AND2X4 U220 ( .A(\mul_a2/fa1_s0_r[24] ), .B(\mul_a2/fa1_s1_r[24] ), 
        .Z(n221) );
  HS65_GSS_XOR2X3 U221 ( .A(\mul_a2/fa1_s0_r[25] ), .B(\mul_a2/fa1_s1_r[25] ), 
        .Z(n236) );
  HS65_GS_NAND2X2 U222 ( .A(n237), .B(n236), .Z(n235) );
  HS65_GS_IVX2 U223 ( .A(n235), .Z(n223) );
  HS65_GS_FA1X4 U224 ( .A0(\mul_a2/fa1_s2_r[25] ), .B0(\mul_a2/fa1_c1_r[24] ), 
        .CI(n221), .CO(n222), .S0(n237) );
  HS65_GS_AOI12X2 U225 ( .A(n236), .B(n237), .C(n222), .Z(n225) );
  HS65_GS_AOI13X2 U226 ( .A(n223), .B(\mul_a2/fa1_c1_r[24] ), .C(
        \mul_a2/fa1_s2_r[25] ), .D(n225), .Z(n385) );
  HS65_GS_AND2X4 U227 ( .A(\mul_a2/fa1_s1_r[25] ), .B(\mul_a2/fa1_s0_r[25] ), 
        .Z(n387) );
  HS65_GS_NAND2X2 U228 ( .A(n224), .B(\mul_a2/fa1_s0_r[26] ), .Z(n386) );
  HS65_GS_OAI21X2 U229 ( .A(n224), .B(\mul_a2/fa1_s0_r[26] ), .C(n386), .Z(
        n384) );
  HS65_GS_AO12X4 U230 ( .A(n385), .B(n384), .C(n225), .Z(n1696) );
  HS65_GS_AND2X4 U231 ( .A(\mul_a2/fa1_s0_r[22] ), .B(\mul_a2/fa1_s1_r[22] ), 
        .Z(n226) );
  HS65_GSS_XOR2X3 U232 ( .A(\mul_a2/fa1_s0_r[23] ), .B(\mul_a2/fa1_s1_r[23] ), 
        .Z(n244) );
  HS65_GS_NAND2X2 U233 ( .A(n245), .B(n244), .Z(n243) );
  HS65_GS_IVX2 U234 ( .A(n243), .Z(n228) );
  HS65_GS_FA1X4 U235 ( .A0(\mul_a2/fa1_s2_r[23] ), .B0(\mul_a2/fa1_c1_r[22] ), 
        .CI(n226), .CO(n227), .S0(n245) );
  HS65_GS_NOR2X2 U236 ( .A(n228), .B(n227), .Z(n229) );
  HS65_GS_AOI13X2 U237 ( .A(n228), .B(\mul_a2/fa1_s2_r[23] ), .C(
        \mul_a2/fa1_c1_r[22] ), .D(n229), .Z(n380) );
  HS65_GS_AND2X4 U238 ( .A(\mul_a2/fa1_s0_r[23] ), .B(\mul_a2/fa1_s1_r[23] ), 
        .Z(n231) );
  HS65_GSS_XOR2X3 U239 ( .A(\mul_a2/fa1_s0_r[24] ), .B(\mul_a2/fa1_s1_r[24] ), 
        .Z(n233) );
  HS65_GS_NAND2X2 U240 ( .A(n232), .B(n233), .Z(n230) );
  HS65_GS_OAI21X2 U241 ( .A(n232), .B(n233), .C(n230), .Z(n379) );
  HS65_GS_NAND2X2 U242 ( .A(n380), .B(n379), .Z(n378) );
  HS65_GS_NOR2AX3 U243 ( .A(n378), .B(n229), .Z(n1214) );
  HS65_GS_IVX2 U244 ( .A(n230), .Z(n383) );
  HS65_GS_FA1X4 U245 ( .A0(\mul_a2/fa1_s2_r[24] ), .B0(\mul_a2/fa1_c1_r[23] ), 
        .CI(n231), .CO(n382), .S0(n232) );
  HS65_GS_AOI12X2 U246 ( .A(n233), .B(n232), .C(n382), .Z(n234) );
  HS65_GS_AOI13X2 U247 ( .A(n383), .B(\mul_a2/fa1_c1_r[23] ), .C(
        \mul_a2/fa1_s2_r[24] ), .D(n234), .Z(n239) );
  HS65_GS_OAI21X2 U248 ( .A(n237), .B(n236), .C(n235), .Z(n238) );
  HS65_GS_NAND2X2 U249 ( .A(n239), .B(n238), .Z(n381) );
  HS65_GS_OAI21X2 U250 ( .A(n239), .B(n238), .C(n381), .Z(n1213) );
  HS65_GS_AND2X4 U251 ( .A(\mul_a2/fa1_s0_r[21] ), .B(\mul_a2/fa1_s1_r[21] ), 
        .Z(n240) );
  HS65_GSS_XOR2X3 U252 ( .A(\mul_a2/fa1_s0_r[22] ), .B(\mul_a2/fa1_s1_r[22] ), 
        .Z(n252) );
  HS65_GS_NAND2X2 U253 ( .A(n253), .B(n252), .Z(n251) );
  HS65_GS_IVX2 U254 ( .A(n251), .Z(n242) );
  HS65_GS_FA1X4 U255 ( .A0(\mul_a2/fa1_s2_r[22] ), .B0(\mul_a2/fa1_c1_r[21] ), 
        .CI(n240), .CO(n241), .S0(n253) );
  HS65_GS_AOI12X2 U256 ( .A(n252), .B(n253), .C(n241), .Z(n246) );
  HS65_GS_AOI13X2 U257 ( .A(n242), .B(\mul_a2/fa1_c1_r[21] ), .C(
        \mul_a2/fa1_s2_r[22] ), .D(n246), .Z(n248) );
  HS65_GS_OAI21X2 U258 ( .A(n245), .B(n244), .C(n243), .Z(n247) );
  HS65_GS_AOI12X2 U259 ( .A(n248), .B(n247), .C(n246), .Z(n1210) );
  HS65_GSS_XOR2X3 U260 ( .A(n248), .B(n247), .Z(n914) );
  HS65_GS_AND2X4 U261 ( .A(\mul_a2/fa1_s0_r[20] ), .B(\mul_a2/fa1_s1_r[20] ), 
        .Z(n249) );
  HS65_GSS_XOR2X3 U262 ( .A(\mul_a2/fa1_s0_r[21] ), .B(\mul_a2/fa1_s1_r[21] ), 
        .Z(n368) );
  HS65_GS_NAND2X2 U263 ( .A(n369), .B(n368), .Z(n367) );
  HS65_GS_IVX2 U264 ( .A(n367), .Z(n256) );
  HS65_GS_FA1X4 U265 ( .A0(\mul_a2/fa1_s2_r[21] ), .B0(\mul_a2/fa1_c1_r[20] ), 
        .CI(n249), .CO(n255), .S0(n369) );
  HS65_GS_AOI12X2 U266 ( .A(n368), .B(n369), .C(n255), .Z(n250) );
  HS65_GS_AOI13X2 U267 ( .A(n256), .B(\mul_a2/fa1_c1_r[20] ), .C(
        \mul_a2/fa1_s2_r[21] ), .D(n250), .Z(n372) );
  HS65_GS_OAI21X2 U268 ( .A(n253), .B(n252), .C(n251), .Z(n371) );
  HS65_GS_NAND2X2 U269 ( .A(n372), .B(n371), .Z(n254) );
  HS65_GS_OAI21X2 U270 ( .A(n256), .B(n255), .C(n254), .Z(n911) );
  HS65_GSS_XOR2X3 U271 ( .A(\mul_a2/fa1_s0_r[19] ), .B(\mul_a2/fa1_s1_r[19] ), 
        .Z(n266) );
  HS65_GS_AND2X4 U272 ( .A(\mul_a2/fa1_s0_r[18] ), .B(\mul_a2/fa1_s1_r[18] ), 
        .Z(n257) );
  HS65_GS_FA1X4 U273 ( .A0(\mul_a2/fa1_s2_r[19] ), .B0(\mul_a2/fa1_c1_r[18] ), 
        .CI(n257), .CO(n258), .S0(n267) );
  HS65_GS_AOI12X2 U274 ( .A(n266), .B(n267), .C(n258), .Z(n261) );
  HS65_GS_NAND2X2 U275 ( .A(n267), .B(n266), .Z(n265) );
  HS65_GS_IVX2 U276 ( .A(n265), .Z(n259) );
  HS65_GS_AOI13X2 U277 ( .A(n259), .B(\mul_a2/fa1_c1_r[18] ), .C(
        \mul_a2/fa1_s2_r[19] ), .D(n261), .Z(n360) );
  HS65_GS_AND2X4 U278 ( .A(\mul_a2/fa1_s1_r[19] ), .B(\mul_a2/fa1_s0_r[19] ), 
        .Z(n363) );
  HS65_GSS_XOR2X3 U279 ( .A(\mul_a2/fa1_s0_r[20] ), .B(\mul_a2/fa1_s1_r[20] ), 
        .Z(n365) );
  HS65_GS_NAND2X2 U280 ( .A(n364), .B(n365), .Z(n362) );
  HS65_GS_OAI21X2 U281 ( .A(n364), .B(n365), .C(n362), .Z(n359) );
  HS65_GS_AND2X4 U282 ( .A(n360), .B(n359), .Z(n260) );
  HS65_GS_NOR2X2 U283 ( .A(n261), .B(n260), .Z(n902) );
  HS65_GSS_XOR2X3 U284 ( .A(\mul_a2/fa1_s0_r[18] ), .B(\mul_a2/fa1_s1_r[18] ), 
        .Z(n350) );
  HS65_GS_FA1X4 U285 ( .A0(\mul_a2/fa1_s2_r[18] ), .B0(\mul_a2/fa1_c1_r[17] ), 
        .CI(n262), .CO(n263), .S0(n351) );
  HS65_GS_AOI12X2 U286 ( .A(n350), .B(n351), .C(n263), .Z(n269) );
  HS65_GS_NAND2X2 U287 ( .A(n351), .B(n350), .Z(n349) );
  HS65_GS_IVX2 U288 ( .A(n349), .Z(n264) );
  HS65_GS_AOI13X2 U289 ( .A(n264), .B(\mul_a2/fa1_c1_r[17] ), .C(
        \mul_a2/fa1_s2_r[18] ), .D(n269), .Z(n271) );
  HS65_GS_OAI21X2 U290 ( .A(n267), .B(n266), .C(n265), .Z(n270) );
  HS65_GS_AND2X4 U291 ( .A(n271), .B(n270), .Z(n268) );
  HS65_GS_NOR2X2 U292 ( .A(n269), .B(n268), .Z(n357) );
  HS65_GSS_XOR2X3 U293 ( .A(n271), .B(n270), .Z(n899) );
  HS65_GS_FA1X4 U294 ( .A0(\mul_a2/fa1_s2_r[16] ), .B0(\mul_a2/fa1_c1_r[15] ), 
        .CI(n272), .CO(n273), .S0(n281) );
  HS65_GS_AOI12X2 U295 ( .A(n280), .B(n281), .C(n273), .Z(n276) );
  HS65_GS_NAND2X2 U296 ( .A(n281), .B(n280), .Z(n279) );
  HS65_GS_IVX2 U297 ( .A(n279), .Z(n274) );
  HS65_GS_AOI13X2 U298 ( .A(n274), .B(\mul_a2/fa1_c1_r[15] ), .C(
        \mul_a2/fa1_s2_r[16] ), .D(n276), .Z(n342) );
  HS65_GS_FA1X4 U299 ( .A0(\mul_a2/fa1_s0_r[16] ), .B0(\mul_a2/fa1_s1_r[16] ), 
        .CI(\mul_a2/fa1_c0_r[15] ), .CO(n345), .S0(n280) );
  HS65_GS_FA1X4 U300 ( .A0(\mul_a2/fa1_s0_r[17] ), .B0(\mul_a2/fa1_s1_r[17] ), 
        .CI(\mul_a2/fa1_c0_r[16] ), .CO(n262), .S0(n347) );
  HS65_GS_NAND2X2 U301 ( .A(n346), .B(n347), .Z(n344) );
  HS65_GS_OAI21X2 U302 ( .A(n346), .B(n347), .C(n344), .Z(n341) );
  HS65_GS_AND2X4 U303 ( .A(n342), .B(n341), .Z(n275) );
  HS65_GS_NOR2X2 U304 ( .A(n276), .B(n275), .Z(n1200) );
  HS65_GSS_XOR2X3 U305 ( .A(\mul_a2/fa1_c1_r[14] ), .B(\mul_a2/fa1_s2_r[15] ), 
        .Z(n288) );
  HS65_GS_FA1X4 U306 ( .A0(\mul_a2/fa1_s0_r[15] ), .B0(\mul_a2/fa1_s1_r[15] ), 
        .CI(\mul_a2/fa1_c0_r[14] ), .CO(n272), .S0(n287) );
  HS65_GS_AOI12X2 U307 ( .A(\mul_a2/fa1_s2_r[15] ), .B(\mul_a2/fa1_c1_r[14] ), 
        .C(n277), .Z(n283) );
  HS65_GS_AND2X4 U308 ( .A(\mul_a2/fa1_c1_r[14] ), .B(\mul_a2/fa1_s2_r[15] ), 
        .Z(n278) );
  HS65_GS_AOI13X2 U309 ( .A(n278), .B(n286), .C(n287), .D(n283), .Z(n285) );
  HS65_GS_OAI21X2 U310 ( .A(n281), .B(n280), .C(n279), .Z(n284) );
  HS65_GS_AND2X4 U311 ( .A(n285), .B(n284), .Z(n282) );
  HS65_GS_NOR2X2 U312 ( .A(n283), .B(n282), .Z(n339) );
  HS65_GSS_XOR2X3 U313 ( .A(n285), .B(n284), .Z(n894) );
  HS65_GS_FA1X4 U314 ( .A0(n288), .B0(n287), .CI(n286), .CO(n277), .S0(n291)
         );
  HS65_GS_AND2X4 U315 ( .A(\mul_a2/fa1_c1_r[13] ), .B(\mul_a2/fa1_s2_r[14] ), 
        .Z(n290) );
  HS65_GSS_XOR2X3 U316 ( .A(\mul_a2/fa1_c1_r[13] ), .B(\mul_a2/fa1_s2_r[14] ), 
        .Z(n294) );
  HS65_GS_FA1X4 U317 ( .A0(\mul_a2/fa1_s0_r[14] ), .B0(\mul_a2/fa1_s1_r[14] ), 
        .CI(\mul_a2/fa1_c0_r[13] ), .CO(n286), .S0(n293) );
  HS65_GS_IVX2 U318 ( .A(n873), .Z(n874) );
  HS65_GS_FA1X4 U319 ( .A0(n291), .B0(n290), .CI(n289), .CO(n873), .S0(n1193)
         );
  HS65_GS_FA1X4 U320 ( .A0(n294), .B0(n293), .CI(n292), .CO(n289), .S0(n337)
         );
  HS65_GS_FA1X4 U321 ( .A0(\mul_a2/fa1_s0_r[13] ), .B0(\mul_a2/fa1_s1_r[13] ), 
        .CI(\mul_a2/fa1_c0_r[12] ), .CO(n292), .S0(n329) );
  HS65_GS_NAND2X2 U322 ( .A(n337), .B(n336), .Z(n338) );
  HS65_GS_FA1X4 U323 ( .A0(\mul_a2/fa1_s0_r[11] ), .B0(\mul_a2/fa1_s1_r[11] ), 
        .CI(\mul_a2/fa1_c0_r[10] ), .CO(n332), .S0(n321) );
  HS65_GS_FA1X4 U324 ( .A0(\mul_a2/fa1_s0_r[12] ), .B0(\mul_a2/fa1_s1_r[12] ), 
        .CI(\mul_a2/fa1_c0_r[11] ), .CO(n330), .S0(n331) );
  HS65_GS_AND2X4 U325 ( .A(\mul_a2/fa1_s0_r[8] ), .B(\mul_a2/fa1_c0_r[7] ), 
        .Z(n295) );
  HS65_GS_AND2X4 U326 ( .A(n295), .B(n313), .Z(n318) );
  HS65_GS_FA1X4 U327 ( .A0(\mul_a2/fa1_s0_r[10] ), .B0(\mul_a2/fa1_s1_r[10] ), 
        .CI(\mul_a2/fa1_c0_r[9] ), .CO(n322), .S0(n319) );
  HS65_GS_FA1X4 U328 ( .A0(\mul_a2/fa1_s0_r[9] ), .B0(\mul_a2/fa1_s1_r[9] ), 
        .CI(\mul_a2/fa1_c0_r[8] ), .CO(n320), .S0(n313) );
  HS65_GSS_XOR2X3 U329 ( .A(n319), .B(n320), .Z(n317) );
  HS65_GS_AND2X4 U330 ( .A(\mul_a2/fa1_s0_r[6] ), .B(\mul_a2/fa1_c0_r[5] ), 
        .Z(n296) );
  HS65_GSS_XOR2X3 U331 ( .A(\mul_a2/fa1_c0_r[6] ), .B(\mul_a2/fa1_s0_r[7] ), 
        .Z(n306) );
  HS65_GS_AND2X4 U332 ( .A(n296), .B(n306), .Z(n310) );
  HS65_GSS_XOR2X3 U333 ( .A(\mul_a2/fa1_c0_r[7] ), .B(\mul_a2/fa1_s0_r[8] ), 
        .Z(n312) );
  HS65_GS_AND2X4 U334 ( .A(\mul_a2/fa1_s0_r[4] ), .B(\mul_a2/fa1_c0_r[3] ), 
        .Z(n297) );
  HS65_GSS_XOR2X3 U335 ( .A(\mul_a2/fa1_c0_r[4] ), .B(\mul_a2/fa1_s0_r[5] ), 
        .Z(n301) );
  HS65_GS_AND2X4 U336 ( .A(n297), .B(n301), .Z(n303) );
  HS65_GSS_XOR2X3 U337 ( .A(\mul_a2/fa1_c0_r[5] ), .B(\mul_a2/fa1_s0_r[6] ), 
        .Z(n305) );
  HS65_GS_AND2X4 U338 ( .A(\mul_a2/fa1_c0_r[2] ), .B(\mul_a2/fa1_s0_r[3] ), 
        .Z(n299) );
  HS65_GSS_XOR2X3 U339 ( .A(\mul_a2/fa1_c0_r[3] ), .B(\mul_a2/fa1_s0_r[4] ), 
        .Z(n298) );
  HS65_GS_AND2X4 U340 ( .A(n299), .B(n298), .Z(n300) );
  HS65_GS_AND2X4 U341 ( .A(n301), .B(n300), .Z(n302) );
  HS65_GS_PAO2X4 U342 ( .A(n303), .B(n305), .P(n302), .Z(n308) );
  HS65_GS_AND2X4 U343 ( .A(\mul_a2/fa1_s0_r[5] ), .B(\mul_a2/fa1_c0_r[4] ), 
        .Z(n304) );
  HS65_GS_AND2X4 U344 ( .A(n305), .B(n304), .Z(n307) );
  HS65_GS_PAO2X4 U345 ( .A(n308), .B(n307), .P(n306), .Z(n309) );
  HS65_GS_PAO2X4 U346 ( .A(n310), .B(n312), .P(n309), .Z(n315) );
  HS65_GS_AND2X4 U347 ( .A(\mul_a2/fa1_s0_r[7] ), .B(\mul_a2/fa1_c0_r[6] ), 
        .Z(n311) );
  HS65_GS_AND2X4 U348 ( .A(n312), .B(n311), .Z(n314) );
  HS65_GS_PAO2X4 U349 ( .A(n315), .B(n314), .P(n313), .Z(n316) );
  HS65_GS_PAO2X4 U350 ( .A(n318), .B(n317), .P(n316), .Z(n325) );
  HS65_GS_AND2X4 U351 ( .A(n320), .B(n319), .Z(n324) );
  HS65_GS_FA1X4 U352 ( .A0(\mul_a2/fa1_c1_r[10] ), .B0(n322), .CI(n321), .CO(
        n328), .S0(n323) );
  HS65_GS_PAO2X4 U353 ( .A(n325), .B(n324), .P(n323), .Z(n326) );
  HS65_GS_PAO2X4 U354 ( .A(n328), .B(n327), .P(n326), .Z(n335) );
  HS65_GS_FA1X4 U355 ( .A0(\mul_a2/fa1_c1_r[12] ), .B0(n330), .CI(n329), .CO(
        n336), .S0(n334) );
  HS65_GS_FA1X4 U356 ( .A0(\mul_a2/fa1_c1_r[11] ), .B0(n332), .CI(n331), .CO(
        n333), .S0(n327) );
  HS65_GS_PAO2X4 U357 ( .A(n335), .B(n334), .P(n333), .Z(n1189) );
  HS65_GSS_XOR2X3 U358 ( .A(n337), .B(n336), .Z(n1188) );
  HS65_GS_NAND2X2 U359 ( .A(n1189), .B(n1188), .Z(n1187) );
  HS65_GS_NAND2X2 U360 ( .A(n338), .B(n1187), .Z(n1192) );
  HS65_GS_NAND2X2 U361 ( .A(n1193), .B(n1192), .Z(n1191) );
  HS65_GS_PAOI2X1 U362 ( .A(n894), .B(n874), .P(n1191), .Z(n340) );
  HS65_GS_NAND2X2 U363 ( .A(n339), .B(n340), .Z(n343) );
  HS65_GSS_XOR2X3 U364 ( .A(n340), .B(n339), .Z(n1197) );
  HS65_GSS_XNOR2X3 U365 ( .A(n342), .B(n341), .Z(n1196) );
  HS65_GS_NAND2X2 U366 ( .A(n1197), .B(n1196), .Z(n1195) );
  HS65_GS_NAND2X2 U367 ( .A(n343), .B(n1195), .Z(n1199) );
  HS65_GS_IVX2 U368 ( .A(n344), .Z(n356) );
  HS65_GS_FA1X4 U369 ( .A0(\mul_a2/fa1_s2_r[17] ), .B0(\mul_a2/fa1_c1_r[16] ), 
        .CI(n345), .CO(n355), .S0(n346) );
  HS65_GS_AOI12X2 U370 ( .A(n347), .B(n346), .C(n355), .Z(n348) );
  HS65_GS_AOI13X2 U371 ( .A(n356), .B(\mul_a2/fa1_c1_r[16] ), .C(
        \mul_a2/fa1_s2_r[17] ), .D(n348), .Z(n353) );
  HS65_GS_OAI21X2 U372 ( .A(n351), .B(n350), .C(n349), .Z(n352) );
  HS65_GSS_XNOR2X3 U373 ( .A(n353), .B(n352), .Z(n1202) );
  HS65_GS_PAOI2X1 U374 ( .A(n1200), .B(n1199), .P(n1202), .Z(n897) );
  HS65_GS_NAND2X2 U375 ( .A(n353), .B(n352), .Z(n354) );
  HS65_GS_OAI21X2 U376 ( .A(n356), .B(n355), .C(n354), .Z(n896) );
  HS65_GS_PAOI2X1 U377 ( .A(n899), .B(n897), .P(n896), .Z(n358) );
  HS65_GS_NAND2X2 U378 ( .A(n357), .B(n358), .Z(n361) );
  HS65_GSS_XOR2X3 U379 ( .A(n358), .B(n357), .Z(n1206) );
  HS65_GSS_XNOR2X3 U380 ( .A(n360), .B(n359), .Z(n1205) );
  HS65_GS_NAND2X2 U381 ( .A(n1206), .B(n1205), .Z(n1204) );
  HS65_GS_NAND2X2 U382 ( .A(n361), .B(n1204), .Z(n901) );
  HS65_GS_IVX2 U383 ( .A(n362), .Z(n377) );
  HS65_GS_FA1X4 U384 ( .A0(\mul_a2/fa1_s2_r[20] ), .B0(\mul_a2/fa1_c1_r[19] ), 
        .CI(n363), .CO(n376), .S0(n364) );
  HS65_GS_AOI12X2 U385 ( .A(n365), .B(n364), .C(n376), .Z(n366) );
  HS65_GS_AOI13X2 U386 ( .A(n377), .B(\mul_a2/fa1_c1_r[19] ), .C(
        \mul_a2/fa1_s2_r[20] ), .D(n366), .Z(n374) );
  HS65_GS_OAI21X2 U387 ( .A(n369), .B(n368), .C(n367), .Z(n373) );
  HS65_GSS_XOR2X3 U388 ( .A(n374), .B(n373), .Z(n904) );
  HS65_GS_IVX2 U389 ( .A(n904), .Z(n370) );
  HS65_GS_PAOI2X1 U390 ( .A(n902), .B(n901), .P(n370), .Z(n907) );
  HS65_GSS_XOR2X3 U391 ( .A(n372), .B(n371), .Z(n909) );
  HS65_GS_NAND2X2 U392 ( .A(n374), .B(n373), .Z(n375) );
  HS65_GS_OAI21X2 U393 ( .A(n377), .B(n376), .C(n375), .Z(n906) );
  HS65_GS_PAO2X4 U394 ( .A(n907), .B(n909), .P(n906), .Z(n912) );
  HS65_GS_PAOI2X1 U395 ( .A(n914), .B(n911), .P(n912), .Z(n1209) );
  HS65_GS_OAI21X2 U396 ( .A(n380), .B(n379), .C(n378), .Z(n1208) );
  HS65_GS_OA12X4 U397 ( .A(n383), .B(n382), .C(n381), .Z(n916) );
  HS65_GSS_XNOR2X3 U398 ( .A(n385), .B(n384), .Z(n918) );
  HS65_GS_PAOI2X1 U399 ( .A(n917), .B(n916), .P(n918), .Z(n1695) );
  HS65_GS_IVX2 U400 ( .A(n386), .Z(n395) );
  HS65_GS_FA1X4 U401 ( .A0(\mul_a2/fa1_s2_r[26] ), .B0(\mul_a2/fa1_c1_r[25] ), 
        .CI(n387), .CO(n394), .S0(n224) );
  HS65_GS_NOR2X2 U402 ( .A(n395), .B(n394), .Z(n388) );
  HS65_GS_AOI13X2 U403 ( .A(n395), .B(\mul_a2/fa1_s2_r[26] ), .C(
        \mul_a2/fa1_c1_r[25] ), .D(n388), .Z(n392) );
  HS65_GS_OAI21X2 U404 ( .A(n390), .B(\mul_a2/fa1_s0_r[27] ), .C(n389), .Z(
        n391) );
  HS65_GS_NAND2X2 U405 ( .A(n392), .B(n391), .Z(n393) );
  HS65_GS_OA12X4 U406 ( .A(n392), .B(n391), .C(n393), .Z(n1694) );
  HS65_GS_OAI21X2 U407 ( .A(n395), .B(n394), .C(n393), .Z(n1699) );
  HS65_GS_OA12X4 U408 ( .A(n398), .B(n397), .C(n396), .Z(n1698) );
  HS65_GS_OA12X4 U409 ( .A(n401), .B(n400), .C(n399), .Z(n878) );
  HS65_GS_AOI12X2 U410 ( .A(\mul_a2/fa1_s0_r[29] ), .B(n403), .C(n402), .Z(
        n404) );
  HS65_GS_IVX2 U411 ( .A(n404), .Z(n405) );
  HS65_GS_MUXI21X2 U412 ( .D0(n407), .D1(n406), .S0(n405), .Z(n875) );
  HS65_GS_AND2X4 U413 ( .A(\mul_a2/fa1_c1_r[29] ), .B(\mul_a2/fa1_s2_r[30] ), 
        .Z(n413) );
  HS65_GSS_XOR2X3 U414 ( .A(n408), .B(\mul_a2/fa1_s0_r[31] ), .Z(n412) );
  HS65_GS_AND2X4 U415 ( .A(\mul_a2/fa1_s0_r[30] ), .B(n409), .Z(n411) );
  HS65_GS_IVX2 U416 ( .A(n410), .Z(n884) );
  HS65_GS_FA1X4 U417 ( .A0(n413), .B0(n412), .CI(n411), .CO(n414), .S0(n410)
         );
  HS65_GS_IVX2 U418 ( .A(n414), .Z(n881) );
  HS65_GSS_XOR2X3 U419 ( .A(n416), .B(n415), .Z(n417) );
  HS65_GSS_XOR3X2 U420 ( .A(n418), .B(\mul_a2/fa1_c1_r[32] ), .C(n417), .Z(
        n420) );
  HS65_GSS_XOR2X3 U421 ( .A(n420), .B(n419), .Z(n421) );
  HS65_GSS_XOR2X3 U422 ( .A(\mul_a2/fa1_s0_r[33] ), .B(n421), .Z(n422) );
  HS65_GSS_XOR2X3 U423 ( .A(\mul_a2/fa1_s2_r[33] ), .B(n422), .Z(
        \mul_a2/result_sat[15] ) );
  HS65_GS_BFX4 U424 ( .A(valid_in), .Z(n1305) );
  HS65_GS_BFX4 U425 ( .A(n1305), .Z(n1714) );
  HS65_GS_AND2X4 U426 ( .A(\mul_b2/fa1_s0_r[31] ), .B(\mul_b2/fa1_s1_r[31] ), 
        .Z(n519) );
  HS65_GS_NAND2X2 U427 ( .A(\mul_b2/fa1_s0_r[32] ), .B(\mul_b2/fa1_s1_r[32] ), 
        .Z(n521) );
  HS65_GS_OA12X4 U428 ( .A(\mul_b2/fa1_s0_r[32] ), .B(\mul_b2/fa1_s1_r[32] ), 
        .C(n521), .Z(n518) );
  HS65_GS_AND2X4 U429 ( .A(\mul_b2/fa1_s0_r[30] ), .B(\mul_b2/fa1_s1_r[30] ), 
        .Z(n424) );
  HS65_GSS_XOR2X3 U430 ( .A(\mul_b2/fa1_s0_r[31] ), .B(\mul_b2/fa1_s1_r[31] ), 
        .Z(n423) );
  HS65_GS_FA1X4 U431 ( .A0(\mul_b2/fa1_s2_r[31] ), .B0(n424), .CI(n423), .CO(
        n941), .S0(n933) );
  HS65_GS_AND2X4 U432 ( .A(\mul_b2/fa1_s0_r[29] ), .B(\mul_b2/fa1_s1_r[29] ), 
        .Z(n426) );
  HS65_GSS_XOR2X3 U433 ( .A(\mul_b2/fa1_s0_r[30] ), .B(\mul_b2/fa1_s1_r[30] ), 
        .Z(n425) );
  HS65_GS_FA1X4 U434 ( .A0(\mul_b2/fa1_s2_r[30] ), .B0(n426), .CI(n425), .CO(
        n932), .S0(n936) );
  HS65_GS_AND2X4 U435 ( .A(\mul_b2/fa1_s0_r[28] ), .B(\mul_b2/fa1_s1_r[28] ), 
        .Z(n428) );
  HS65_GSS_XOR2X3 U436 ( .A(\mul_b2/fa1_s0_r[29] ), .B(\mul_b2/fa1_s1_r[29] ), 
        .Z(n427) );
  HS65_GS_FA1X4 U437 ( .A0(\mul_b2/fa1_s2_r[29] ), .B0(n428), .CI(n427), .CO(
        n935), .S0(n939) );
  HS65_GS_AND2X4 U438 ( .A(\mul_b2/fa1_s0_r[27] ), .B(\mul_b2/fa1_s1_r[27] ), 
        .Z(n430) );
  HS65_GSS_XOR2X3 U439 ( .A(\mul_b2/fa1_s0_r[28] ), .B(\mul_b2/fa1_s1_r[28] ), 
        .Z(n429) );
  HS65_GS_FA1X4 U440 ( .A0(\mul_b2/fa1_s2_r[28] ), .B0(n430), .CI(n429), .CO(
        n938), .S0(n1403) );
  HS65_GS_AND2X4 U441 ( .A(\mul_b2/fa1_s0_r[26] ), .B(\mul_b2/fa1_s1_r[26] ), 
        .Z(n512) );
  HS65_GSS_XOR2X3 U442 ( .A(\mul_b2/fa1_s0_r[27] ), .B(\mul_b2/fa1_s1_r[27] ), 
        .Z(n511) );
  HS65_GS_AND2X4 U443 ( .A(\mul_b2/fa1_s0_r[24] ), .B(\mul_b2/fa1_s1_r[24] ), 
        .Z(n432) );
  HS65_GSS_XOR2X3 U444 ( .A(\mul_b2/fa1_s0_r[25] ), .B(\mul_b2/fa1_s1_r[25] ), 
        .Z(n431) );
  HS65_GS_AND2X4 U445 ( .A(\mul_b2/fa1_s0_r[25] ), .B(\mul_b2/fa1_s1_r[25] ), 
        .Z(n514) );
  HS65_GSS_XOR2X3 U446 ( .A(\mul_b2/fa1_s0_r[26] ), .B(\mul_b2/fa1_s1_r[26] ), 
        .Z(n513) );
  HS65_GS_AND2X4 U447 ( .A(\mul_b2/fa1_s0_r[23] ), .B(\mul_b2/fa1_s1_r[23] ), 
        .Z(n434) );
  HS65_GSS_XOR2X3 U448 ( .A(\mul_b2/fa1_s0_r[24] ), .B(\mul_b2/fa1_s1_r[24] ), 
        .Z(n433) );
  HS65_GS_FA1X4 U449 ( .A0(\mul_b2/fa1_s2_r[25] ), .B0(n432), .CI(n431), .CO(
        n510), .S0(n506) );
  HS65_GS_AND2X4 U450 ( .A(\mul_b2/fa1_s0_r[22] ), .B(\mul_b2/fa1_s1_r[22] ), 
        .Z(n436) );
  HS65_GSS_XOR2X3 U451 ( .A(\mul_b2/fa1_s0_r[23] ), .B(\mul_b2/fa1_s1_r[23] ), 
        .Z(n435) );
  HS65_GS_FA1X4 U452 ( .A0(\mul_b2/fa1_s2_r[24] ), .B0(n434), .CI(n433), .CO(
        n507), .S0(n503) );
  HS65_GS_AND2X4 U453 ( .A(\mul_b2/fa1_s0_r[21] ), .B(\mul_b2/fa1_s1_r[21] ), 
        .Z(n438) );
  HS65_GSS_XOR2X3 U454 ( .A(\mul_b2/fa1_s0_r[22] ), .B(\mul_b2/fa1_s1_r[22] ), 
        .Z(n437) );
  HS65_GS_FA1X4 U455 ( .A0(\mul_b2/fa1_s2_r[23] ), .B0(n436), .CI(n435), .CO(
        n504), .S0(n500) );
  HS65_GS_AND2X4 U456 ( .A(\mul_b2/fa1_s0_r[20] ), .B(\mul_b2/fa1_s1_r[20] ), 
        .Z(n440) );
  HS65_GSS_XOR2X3 U457 ( .A(\mul_b2/fa1_s0_r[21] ), .B(\mul_b2/fa1_s1_r[21] ), 
        .Z(n439) );
  HS65_GS_FA1X4 U458 ( .A0(\mul_b2/fa1_s2_r[22] ), .B0(n438), .CI(n437), .CO(
        n501), .S0(n497) );
  HS65_GS_AND2X4 U459 ( .A(\mul_b2/fa1_s0_r[19] ), .B(\mul_b2/fa1_s1_r[19] ), 
        .Z(n442) );
  HS65_GSS_XOR2X3 U460 ( .A(\mul_b2/fa1_s0_r[20] ), .B(\mul_b2/fa1_s1_r[20] ), 
        .Z(n441) );
  HS65_GS_FA1X4 U461 ( .A0(\mul_b2/fa1_s2_r[21] ), .B0(n440), .CI(n439), .CO(
        n498), .S0(n494) );
  HS65_GS_AND2X4 U462 ( .A(\mul_b2/fa1_s0_r[18] ), .B(\mul_b2/fa1_s1_r[18] ), 
        .Z(n444) );
  HS65_GSS_XOR2X3 U463 ( .A(\mul_b2/fa1_s0_r[19] ), .B(\mul_b2/fa1_s1_r[19] ), 
        .Z(n443) );
  HS65_GS_FA1X4 U464 ( .A0(\mul_b2/fa1_s2_r[20] ), .B0(n442), .CI(n441), .CO(
        n495), .S0(n491) );
  HS65_GS_AND2X4 U465 ( .A(\mul_b2/fa1_s0_r[17] ), .B(\mul_b2/fa1_s1_r[17] ), 
        .Z(n446) );
  HS65_GSS_XOR2X3 U466 ( .A(\mul_b2/fa1_s0_r[18] ), .B(\mul_b2/fa1_s1_r[18] ), 
        .Z(n445) );
  HS65_GS_FA1X4 U467 ( .A0(\mul_b2/fa1_s2_r[19] ), .B0(n444), .CI(n443), .CO(
        n492), .S0(n488) );
  HS65_GS_AND2X4 U468 ( .A(\mul_b2/fa1_s0_r[16] ), .B(\mul_b2/fa1_s1_r[16] ), 
        .Z(n448) );
  HS65_GSS_XOR2X3 U469 ( .A(\mul_b2/fa1_s0_r[17] ), .B(\mul_b2/fa1_s1_r[17] ), 
        .Z(n447) );
  HS65_GS_FA1X4 U470 ( .A0(\mul_b2/fa1_s2_r[18] ), .B0(n446), .CI(n445), .CO(
        n489), .S0(n485) );
  HS65_GS_AND2X4 U471 ( .A(\mul_b2/fa1_s0_r[15] ), .B(\mul_b2/fa1_s1_r[15] ), 
        .Z(n450) );
  HS65_GSS_XOR2X3 U472 ( .A(\mul_b2/fa1_s0_r[16] ), .B(\mul_b2/fa1_s1_r[16] ), 
        .Z(n449) );
  HS65_GS_FA1X4 U473 ( .A0(\mul_b2/fa1_s2_r[17] ), .B0(n448), .CI(n447), .CO(
        n486), .S0(n482) );
  HS65_GS_AND2X4 U474 ( .A(\mul_b2/fa1_s0_r[14] ), .B(\mul_b2/fa1_s1_r[14] ), 
        .Z(n453) );
  HS65_GSS_XOR2X3 U475 ( .A(\mul_b2/fa1_s0_r[15] ), .B(\mul_b2/fa1_s1_r[15] ), 
        .Z(n452) );
  HS65_GS_FA1X4 U476 ( .A0(\mul_b2/fa1_s2_r[16] ), .B0(n450), .CI(n449), .CO(
        n483), .S0(n479) );
  HS65_GS_NOR2X2 U477 ( .A(n480), .B(n479), .Z(n451) );
  HS65_GS_AOI12X2 U478 ( .A(n479), .B(n480), .C(n451), .Z(n960) );
  HS65_GS_AND2X4 U479 ( .A(\mul_b2/fa1_s0_r[13] ), .B(\mul_b2/fa1_s1_r[13] ), 
        .Z(n455) );
  HS65_GSS_XOR2X3 U480 ( .A(\mul_b2/fa1_s0_r[14] ), .B(\mul_b2/fa1_s1_r[14] ), 
        .Z(n454) );
  HS65_GS_FA1X4 U481 ( .A0(\mul_b2/fa1_s2_r[15] ), .B0(n453), .CI(n452), .CO(
        n480), .S0(n476) );
  HS65_GS_NAND2X2 U482 ( .A(\mul_b2/fa1_s0_r[12] ), .B(\mul_b2/fa1_s1_r[12] ), 
        .Z(n458) );
  HS65_GS_IVX2 U483 ( .A(n458), .Z(n457) );
  HS65_GSS_XOR2X3 U484 ( .A(\mul_b2/fa1_s0_r[13] ), .B(\mul_b2/fa1_s1_r[13] ), 
        .Z(n456) );
  HS65_GS_FA1X4 U485 ( .A0(\mul_b2/fa1_s2_r[14] ), .B0(n455), .CI(n454), .CO(
        n477), .S0(n473) );
  HS65_GS_FA1X4 U486 ( .A0(\mul_b2/fa1_s2_r[13] ), .B0(n457), .CI(n456), .CO(
        n474), .S0(n471) );
  HS65_GS_OAI21X2 U487 ( .A(\mul_b2/fa1_s0_r[12] ), .B(\mul_b2/fa1_s1_r[12] ), 
        .C(n458), .Z(n461) );
  HS65_GS_IVX2 U488 ( .A(\mul_b2/fa1_s2_r[12] ), .Z(n460) );
  HS65_GS_NAND2X2 U489 ( .A(\mul_b2/fa1_s1_r[11] ), .B(\mul_b2/fa1_s0_r[11] ), 
        .Z(n459) );
  HS65_GS_PAOI2X1 U490 ( .A(n461), .B(n460), .P(n459), .Z(n470) );
  HS65_GS_AND2X4 U491 ( .A(n461), .B(n460), .Z(n468) );
  HS65_GS_OAI21X2 U492 ( .A(\mul_b2/fa1_s1_r[11] ), .B(\mul_b2/fa1_s0_r[11] ), 
        .C(n471), .Z(n467) );
  HS65_GS_AND2X4 U493 ( .A(\mul_b2/fa1_s0_r[6] ), .B(\mul_b2/fa1_s1_r[6] ), 
        .Z(n462) );
  HS65_GS_PAO2X4 U494 ( .A(\mul_b2/fa1_s0_r[7] ), .B(\mul_b2/fa1_s1_r[7] ), 
        .P(n462), .Z(n463) );
  HS65_GS_PAO2X4 U495 ( .A(\mul_b2/fa1_s1_r[8] ), .B(\mul_b2/fa1_s0_r[8] ), 
        .P(n463), .Z(n464) );
  HS65_GS_PAO2X4 U496 ( .A(\mul_b2/fa1_s1_r[9] ), .B(\mul_b2/fa1_s0_r[9] ), 
        .P(n464), .Z(n465) );
  HS65_GS_PAOI2X1 U497 ( .A(\mul_b2/fa1_s1_r[10] ), .B(\mul_b2/fa1_s0_r[10] ), 
        .P(n465), .Z(n466) );
  HS65_GS_NOR3X1 U498 ( .A(n468), .B(n467), .C(n466), .Z(n469) );
  HS65_GS_AOI12X2 U499 ( .A(n471), .B(n470), .C(n469), .Z(n952) );
  HS65_GS_NAND2X2 U500 ( .A(n473), .B(n474), .Z(n472) );
  HS65_GS_OAI21X2 U501 ( .A(n473), .B(n474), .C(n472), .Z(n951) );
  HS65_GS_NOR2X2 U502 ( .A(n952), .B(n951), .Z(n950) );
  HS65_GS_AOI12X2 U503 ( .A(n474), .B(n473), .C(n950), .Z(n956) );
  HS65_GS_NAND2X2 U504 ( .A(n476), .B(n477), .Z(n475) );
  HS65_GS_OAI21X2 U505 ( .A(n476), .B(n477), .C(n475), .Z(n955) );
  HS65_GS_NOR2X2 U506 ( .A(n956), .B(n955), .Z(n954) );
  HS65_GS_AOI12X2 U507 ( .A(n477), .B(n476), .C(n954), .Z(n959) );
  HS65_GS_NAND2X2 U508 ( .A(n960), .B(n959), .Z(n478) );
  HS65_GS_OAI21X2 U509 ( .A(n480), .B(n479), .C(n478), .Z(n963) );
  HS65_GS_NAND2X2 U510 ( .A(n482), .B(n483), .Z(n481) );
  HS65_GS_OAI21X2 U511 ( .A(n482), .B(n483), .C(n481), .Z(n962) );
  HS65_GS_NOR2X2 U512 ( .A(n963), .B(n962), .Z(n961) );
  HS65_GS_AOI12X2 U513 ( .A(n483), .B(n482), .C(n961), .Z(n967) );
  HS65_GS_NAND2X2 U514 ( .A(n485), .B(n486), .Z(n484) );
  HS65_GS_OAI21X2 U515 ( .A(n485), .B(n486), .C(n484), .Z(n966) );
  HS65_GS_NOR2X2 U516 ( .A(n967), .B(n966), .Z(n965) );
  HS65_GS_AOI12X2 U517 ( .A(n486), .B(n485), .C(n965), .Z(n971) );
  HS65_GS_NAND2X2 U518 ( .A(n488), .B(n489), .Z(n487) );
  HS65_GS_OAI21X2 U519 ( .A(n488), .B(n489), .C(n487), .Z(n970) );
  HS65_GS_NOR2X2 U520 ( .A(n971), .B(n970), .Z(n969) );
  HS65_GS_AOI12X2 U521 ( .A(n489), .B(n488), .C(n969), .Z(n975) );
  HS65_GS_NAND2X2 U522 ( .A(n491), .B(n492), .Z(n490) );
  HS65_GS_OAI21X2 U523 ( .A(n491), .B(n492), .C(n490), .Z(n974) );
  HS65_GS_NOR2X2 U524 ( .A(n975), .B(n974), .Z(n973) );
  HS65_GS_AOI12X2 U525 ( .A(n492), .B(n491), .C(n973), .Z(n979) );
  HS65_GS_NAND2X2 U526 ( .A(n494), .B(n495), .Z(n493) );
  HS65_GS_OAI21X2 U527 ( .A(n494), .B(n495), .C(n493), .Z(n978) );
  HS65_GS_NOR2X2 U528 ( .A(n979), .B(n978), .Z(n977) );
  HS65_GS_AOI12X2 U529 ( .A(n495), .B(n494), .C(n977), .Z(n983) );
  HS65_GS_NAND2X2 U530 ( .A(n497), .B(n498), .Z(n496) );
  HS65_GS_OAI21X2 U531 ( .A(n497), .B(n498), .C(n496), .Z(n982) );
  HS65_GS_NOR2X2 U532 ( .A(n983), .B(n982), .Z(n981) );
  HS65_GS_AOI12X2 U533 ( .A(n498), .B(n497), .C(n981), .Z(n987) );
  HS65_GS_NAND2X2 U534 ( .A(n500), .B(n501), .Z(n499) );
  HS65_GS_OAI21X2 U535 ( .A(n500), .B(n501), .C(n499), .Z(n986) );
  HS65_GS_NOR2X2 U536 ( .A(n987), .B(n986), .Z(n985) );
  HS65_GS_AOI12X2 U537 ( .A(n501), .B(n500), .C(n985), .Z(n991) );
  HS65_GS_NAND2X2 U538 ( .A(n503), .B(n504), .Z(n502) );
  HS65_GS_OAI21X2 U539 ( .A(n503), .B(n504), .C(n502), .Z(n990) );
  HS65_GS_NOR2X2 U540 ( .A(n991), .B(n990), .Z(n989) );
  HS65_GS_AOI12X2 U541 ( .A(n504), .B(n503), .C(n989), .Z(n995) );
  HS65_GS_NAND2X2 U542 ( .A(n506), .B(n507), .Z(n505) );
  HS65_GS_OAI21X2 U543 ( .A(n506), .B(n507), .C(n505), .Z(n994) );
  HS65_GS_NOR2X2 U544 ( .A(n995), .B(n994), .Z(n993) );
  HS65_GS_AOI12X2 U545 ( .A(n507), .B(n506), .C(n993), .Z(n999) );
  HS65_GS_NAND2X2 U546 ( .A(n509), .B(n510), .Z(n508) );
  HS65_GS_OAI21X2 U547 ( .A(n509), .B(n510), .C(n508), .Z(n998) );
  HS65_GS_NOR2X2 U548 ( .A(n999), .B(n998), .Z(n997) );
  HS65_GS_AOI12X2 U549 ( .A(n510), .B(n509), .C(n997), .Z(n1399) );
  HS65_GS_FA1X4 U550 ( .A0(\mul_b2/fa1_s2_r[27] ), .B0(n512), .CI(n511), .CO(
        n1402), .S0(n516) );
  HS65_GS_FA1X4 U551 ( .A0(\mul_b2/fa1_s2_r[26] ), .B0(n514), .CI(n513), .CO(
        n515), .S0(n509) );
  HS65_GS_NAND2X2 U552 ( .A(n516), .B(n515), .Z(n517) );
  HS65_GS_OAI21X2 U553 ( .A(n516), .B(n515), .C(n517), .Z(n1400) );
  HS65_GS_OAI21X2 U554 ( .A(n1399), .B(n1400), .C(n517), .Z(n1401) );
  HS65_GS_FA1X4 U555 ( .A0(\mul_b2/fa1_s2_r[32] ), .B0(n519), .CI(n518), .CO(
        n520), .S0(n942) );
  HS65_GSS_XNOR2X3 U556 ( .A(n521), .B(n520), .Z(n522) );
  HS65_GSS_XOR3X2 U557 ( .A(\mul_b2/fa1_s2_r[33] ), .B(n523), .C(n522), .Z(
        n524) );
  HS65_GSS_XOR3X2 U558 ( .A(\mul_b2/fa1_s1_r[33] ), .B(\mul_b2/fa1_s0_r[33] ), 
        .C(n524), .Z(\mul_b2/result_sat[15] ) );
  HS65_GS_NAND2X2 U559 ( .A(\mul_a1/fa1_s1_r[32] ), .B(\mul_a1/fa1_s0_r[32] ), 
        .Z(n527) );
  HS65_GS_IVX2 U560 ( .A(\mul_a1/fa1_c1_r[31] ), .Z(n525) );
  HS65_GS_NAND2X2 U561 ( .A(\mul_a1/fa1_s1_r[31] ), .B(\mul_a1/fa1_s0_r[31] ), 
        .Z(n529) );
  HS65_GS_OAI21X2 U562 ( .A(\mul_a1/fa1_s1_r[32] ), .B(\mul_a1/fa1_s0_r[32] ), 
        .C(n527), .Z(n528) );
  HS65_GS_PAOI2X1 U563 ( .A(n525), .B(n529), .P(n528), .Z(n526) );
  HS65_GSS_XOR3X2 U564 ( .A(\mul_a1/fa1_s0_r[33] ), .B(n527), .C(n526), .Z(
        n625) );
  HS65_GSS_XOR3X2 U565 ( .A(\mul_a1/fa1_c1_r[31] ), .B(n529), .C(n528), .Z(
        n531) );
  HS65_GS_AND2X4 U566 ( .A(\mul_a1/fa1_s0_r[30] ), .B(\mul_a1/fa1_s1_r[30] ), 
        .Z(n533) );
  HS65_GSS_XOR2X3 U567 ( .A(\mul_a1/fa1_s1_r[31] ), .B(\mul_a1/fa1_s0_r[31] ), 
        .Z(n532) );
  HS65_GS_NAND2X2 U568 ( .A(n531), .B(n530), .Z(n624) );
  HS65_GS_OAI21X2 U569 ( .A(n531), .B(n530), .C(n624), .Z(n1004) );
  HS65_GS_FA1X4 U570 ( .A0(\mul_a1/fa1_c1_r[30] ), .B0(n533), .CI(n532), .CO(
        n530), .S0(n1007) );
  HS65_GS_AND2X4 U571 ( .A(\mul_a1/fa1_s0_r[29] ), .B(\mul_a1/fa1_s1_r[29] ), 
        .Z(n535) );
  HS65_GSS_XOR2X3 U572 ( .A(\mul_a1/fa1_s0_r[30] ), .B(\mul_a1/fa1_s1_r[30] ), 
        .Z(n534) );
  HS65_GS_FA1X4 U573 ( .A0(\mul_a1/fa1_c1_r[29] ), .B0(n535), .CI(n534), .CO(
        n1006), .S0(n1012) );
  HS65_GS_AND2X4 U574 ( .A(\mul_a1/fa1_s0_r[28] ), .B(\mul_a1/fa1_s1_r[28] ), 
        .Z(n537) );
  HS65_GSS_XOR2X3 U575 ( .A(\mul_a1/fa1_s0_r[29] ), .B(\mul_a1/fa1_s1_r[29] ), 
        .Z(n536) );
  HS65_GS_FA1X4 U576 ( .A0(\mul_a1/fa1_c1_r[28] ), .B0(n537), .CI(n536), .CO(
        n1011), .S0(n1015) );
  HS65_GS_AND2X4 U577 ( .A(\mul_a1/fa1_s0_r[27] ), .B(\mul_a1/fa1_s1_r[27] ), 
        .Z(n539) );
  HS65_GSS_XOR2X3 U578 ( .A(\mul_a1/fa1_s0_r[28] ), .B(\mul_a1/fa1_s1_r[28] ), 
        .Z(n538) );
  HS65_GS_FA1X4 U579 ( .A0(\mul_a1/fa1_c1_r[27] ), .B0(n539), .CI(n538), .CO(
        n1014), .S0(n1442) );
  HS65_GS_AND2X4 U580 ( .A(\mul_a1/fa1_s0_r[26] ), .B(\mul_a1/fa1_s1_r[26] ), 
        .Z(n616) );
  HS65_GSS_XOR2X3 U581 ( .A(\mul_a1/fa1_s0_r[27] ), .B(\mul_a1/fa1_s1_r[27] ), 
        .Z(n615) );
  HS65_GS_AND2X4 U582 ( .A(\mul_a1/fa1_s0_r[24] ), .B(\mul_a1/fa1_s1_r[24] ), 
        .Z(n541) );
  HS65_GSS_XOR2X3 U583 ( .A(\mul_a1/fa1_s1_r[25] ), .B(\mul_a1/fa1_s0_r[25] ), 
        .Z(n540) );
  HS65_GS_AND2X4 U584 ( .A(\mul_a1/fa1_s1_r[25] ), .B(\mul_a1/fa1_s0_r[25] ), 
        .Z(n618) );
  HS65_GSS_XOR2X3 U585 ( .A(\mul_a1/fa1_s0_r[26] ), .B(\mul_a1/fa1_s1_r[26] ), 
        .Z(n617) );
  HS65_GS_AND2X4 U586 ( .A(\mul_a1/fa1_s0_r[23] ), .B(\mul_a1/fa1_s1_r[23] ), 
        .Z(n543) );
  HS65_GSS_XOR2X3 U587 ( .A(\mul_a1/fa1_s0_r[24] ), .B(\mul_a1/fa1_s1_r[24] ), 
        .Z(n542) );
  HS65_GS_FA1X4 U588 ( .A0(\mul_a1/fa1_c1_r[24] ), .B0(n541), .CI(n540), .CO(
        n614), .S0(n610) );
  HS65_GS_AND2X4 U589 ( .A(\mul_a1/fa1_s0_r[22] ), .B(\mul_a1/fa1_s1_r[22] ), 
        .Z(n545) );
  HS65_GSS_XOR2X3 U590 ( .A(\mul_a1/fa1_s0_r[23] ), .B(\mul_a1/fa1_s1_r[23] ), 
        .Z(n544) );
  HS65_GS_FA1X4 U591 ( .A0(\mul_a1/fa1_c1_r[23] ), .B0(n543), .CI(n542), .CO(
        n611), .S0(n607) );
  HS65_GS_AND2X4 U592 ( .A(\mul_a1/fa1_s0_r[21] ), .B(\mul_a1/fa1_s1_r[21] ), 
        .Z(n547) );
  HS65_GSS_XOR2X3 U593 ( .A(\mul_a1/fa1_s0_r[22] ), .B(\mul_a1/fa1_s1_r[22] ), 
        .Z(n546) );
  HS65_GS_FA1X4 U594 ( .A0(\mul_a1/fa1_c1_r[22] ), .B0(n545), .CI(n544), .CO(
        n608), .S0(n603) );
  HS65_GS_FA1X4 U595 ( .A0(\mul_a1/fa1_c1_r[21] ), .B0(n547), .CI(n546), .CO(
        n604), .S0(n1027) );
  HS65_GS_AND2X4 U596 ( .A(\mul_a1/fa1_s1_r[20] ), .B(\mul_a1/fa1_s0_r[20] ), 
        .Z(n600) );
  HS65_GSS_XOR2X3 U597 ( .A(\mul_a1/fa1_s0_r[21] ), .B(\mul_a1/fa1_s1_r[21] ), 
        .Z(n599) );
  HS65_GS_AND2X4 U598 ( .A(\mul_a1/fa1_s0_r[15] ), .B(\mul_a1/fa1_s1_r[15] ), 
        .Z(n549) );
  HS65_GSS_XOR2X3 U599 ( .A(\mul_a1/fa1_s1_r[16] ), .B(\mul_a1/fa1_s0_r[16] ), 
        .Z(n548) );
  HS65_GS_AND2X4 U600 ( .A(\mul_a1/fa1_s1_r[16] ), .B(\mul_a1/fa1_s0_r[16] ), 
        .Z(n592) );
  HS65_GSS_XOR2X3 U601 ( .A(\mul_a1/fa1_s1_r[17] ), .B(\mul_a1/fa1_s0_r[17] ), 
        .Z(n591) );
  HS65_GS_AND2X4 U602 ( .A(\mul_a1/fa1_s0_r[14] ), .B(\mul_a1/fa1_s1_r[14] ), 
        .Z(n585) );
  HS65_GSS_XOR2X3 U603 ( .A(\mul_a1/fa1_s0_r[15] ), .B(\mul_a1/fa1_s1_r[15] ), 
        .Z(n584) );
  HS65_GS_FA1X4 U604 ( .A0(\mul_a1/fa1_c1_r[15] ), .B0(n549), .CI(n548), .CO(
        n1418), .S0(n1413) );
  HS65_GS_AND2X4 U605 ( .A(\mul_a1/fa1_s0_r[12] ), .B(\mul_a1/fa1_s1_r[12] ), 
        .Z(n551) );
  HS65_GSS_XOR2X3 U606 ( .A(\mul_a1/fa1_s1_r[13] ), .B(\mul_a1/fa1_s0_r[13] ), 
        .Z(n550) );
  HS65_GS_AND2X4 U607 ( .A(\mul_a1/fa1_s1_r[13] ), .B(\mul_a1/fa1_s0_r[13] ), 
        .Z(n587) );
  HS65_GSS_XOR2X3 U608 ( .A(\mul_a1/fa1_s0_r[14] ), .B(\mul_a1/fa1_s1_r[14] ), 
        .Z(n586) );
  HS65_GS_FA1X4 U609 ( .A0(\mul_a1/fa1_c1_r[12] ), .B0(n551), .CI(n550), .CO(
        n583), .S0(n580) );
  HS65_GS_AND2X4 U610 ( .A(\mul_a1/fa1_s0_r[11] ), .B(\mul_a1/fa1_s1_r[11] ), 
        .Z(n553) );
  HS65_GSS_XOR2X3 U611 ( .A(\mul_a1/fa1_s0_r[12] ), .B(\mul_a1/fa1_s1_r[12] ), 
        .Z(n552) );
  HS65_GS_AND2X4 U612 ( .A(\mul_a1/fa1_s0_r[10] ), .B(\mul_a1/fa1_s1_r[10] ), 
        .Z(n555) );
  HS65_GSS_XOR2X3 U613 ( .A(\mul_a1/fa1_s0_r[11] ), .B(\mul_a1/fa1_s1_r[11] ), 
        .Z(n554) );
  HS65_GS_FA1X4 U614 ( .A0(\mul_a1/fa1_c1_r[11] ), .B0(n553), .CI(n552), .CO(
        n579), .S0(n576) );
  HS65_GS_AND2X4 U615 ( .A(\mul_a1/fa1_s0_r[9] ), .B(\mul_a1/fa1_s1_r[9] ), 
        .Z(n557) );
  HS65_GSS_XOR2X3 U616 ( .A(\mul_a1/fa1_s0_r[10] ), .B(\mul_a1/fa1_s1_r[10] ), 
        .Z(n556) );
  HS65_GS_FA1X4 U617 ( .A0(\mul_a1/fa1_c1_r[10] ), .B0(n555), .CI(n554), .CO(
        n577), .S0(n573) );
  HS65_GS_AND2X4 U618 ( .A(\mul_a1/fa1_s0_r[8] ), .B(\mul_a1/fa1_s1_r[8] ), 
        .Z(n559) );
  HS65_GSS_XOR2X3 U619 ( .A(\mul_a1/fa1_s0_r[9] ), .B(\mul_a1/fa1_s1_r[9] ), 
        .Z(n558) );
  HS65_GS_FA1X4 U620 ( .A0(\mul_a1/fa1_c1_r[9] ), .B0(n557), .CI(n556), .CO(
        n574), .S0(n570) );
  HS65_GS_AND2X4 U621 ( .A(\mul_a1/fa1_s1_r[7] ), .B(\mul_a1/fa1_s0_r[7] ), 
        .Z(n560) );
  HS65_GSS_XOR2X3 U622 ( .A(\mul_a1/fa1_s0_r[8] ), .B(\mul_a1/fa1_s1_r[8] ), 
        .Z(n564) );
  HS65_GS_AND2X4 U623 ( .A(n560), .B(n564), .Z(n568) );
  HS65_GS_FA1X4 U624 ( .A0(\mul_a1/fa1_c1_r[8] ), .B0(n559), .CI(n558), .CO(
        n571), .S0(n567) );
  HS65_GS_NAND2X2 U625 ( .A(\mul_a1/fa1_s0_r[6] ), .B(\mul_a1/fa1_s1_r[6] ), 
        .Z(n563) );
  HS65_GS_IVX2 U626 ( .A(n560), .Z(n561) );
  HS65_GS_OAI21X2 U627 ( .A(\mul_a1/fa1_s1_r[7] ), .B(\mul_a1/fa1_s0_r[7] ), 
        .C(n561), .Z(n562) );
  HS65_GS_NOR2X2 U628 ( .A(n563), .B(n562), .Z(n565) );
  HS65_GS_AND2X4 U629 ( .A(n565), .B(n564), .Z(n566) );
  HS65_GS_PAO2X4 U630 ( .A(n568), .B(n567), .P(n566), .Z(n569) );
  HS65_GS_PAO2X4 U631 ( .A(n571), .B(n570), .P(n569), .Z(n572) );
  HS65_GS_PAO2X4 U632 ( .A(n574), .B(n573), .P(n572), .Z(n575) );
  HS65_GS_PAO2X4 U633 ( .A(n577), .B(n576), .P(n575), .Z(n578) );
  HS65_GS_PAOI2X1 U634 ( .A(n580), .B(n579), .P(n578), .Z(n1024) );
  HS65_GS_NAND2X2 U635 ( .A(n582), .B(n583), .Z(n581) );
  HS65_GS_OAI21X2 U636 ( .A(n582), .B(n583), .C(n581), .Z(n1023) );
  HS65_GS_NOR2X2 U637 ( .A(n1024), .B(n1023), .Z(n1022) );
  HS65_GS_AOI12X2 U638 ( .A(n583), .B(n582), .C(n1022), .Z(n1410) );
  HS65_GS_FA1X4 U639 ( .A0(\mul_a1/fa1_c1_r[14] ), .B0(n585), .CI(n584), .CO(
        n1414), .S0(n589) );
  HS65_GS_FA1X4 U640 ( .A0(\mul_a1/fa1_c1_r[13] ), .B0(n587), .CI(n586), .CO(
        n588), .S0(n582) );
  HS65_GS_NAND2X2 U641 ( .A(n589), .B(n588), .Z(n590) );
  HS65_GS_OAI21X2 U642 ( .A(n589), .B(n588), .C(n590), .Z(n1411) );
  HS65_GS_OAI21X2 U643 ( .A(n1410), .B(n1411), .C(n590), .Z(n1412) );
  HS65_GS_FA1X4 U644 ( .A0(\mul_a1/fa1_c1_r[16] ), .B0(n592), .CI(n591), .CO(
        n1421), .S0(n1417) );
  HS65_GS_AND2X4 U645 ( .A(\mul_a1/fa1_s1_r[17] ), .B(\mul_a1/fa1_s0_r[17] ), 
        .Z(n594) );
  HS65_GSS_XOR2X3 U646 ( .A(\mul_a1/fa1_s1_r[18] ), .B(\mul_a1/fa1_s0_r[18] ), 
        .Z(n593) );
  HS65_GS_FA1X4 U647 ( .A0(\mul_a1/fa1_c1_r[17] ), .B0(n594), .CI(n593), .CO(
        n1425), .S0(n1420) );
  HS65_GS_AND2X4 U648 ( .A(\mul_a1/fa1_s1_r[18] ), .B(\mul_a1/fa1_s0_r[18] ), 
        .Z(n596) );
  HS65_GSS_XOR2X3 U649 ( .A(\mul_a1/fa1_s1_r[19] ), .B(\mul_a1/fa1_s0_r[19] ), 
        .Z(n595) );
  HS65_GS_FA1X4 U650 ( .A0(\mul_a1/fa1_c1_r[18] ), .B0(n596), .CI(n595), .CO(
        n1429), .S0(n1424) );
  HS65_GS_AND2X4 U651 ( .A(\mul_a1/fa1_s1_r[19] ), .B(\mul_a1/fa1_s0_r[19] ), 
        .Z(n598) );
  HS65_GSS_XOR2X3 U652 ( .A(\mul_a1/fa1_s1_r[20] ), .B(\mul_a1/fa1_s0_r[20] ), 
        .Z(n597) );
  HS65_GS_FA1X4 U653 ( .A0(\mul_a1/fa1_c1_r[19] ), .B0(n598), .CI(n597), .CO(
        n1433), .S0(n1428) );
  HS65_GS_FA1X4 U654 ( .A0(\mul_a1/fa1_c1_r[20] ), .B0(n600), .CI(n599), .CO(
        n1026), .S0(n1432) );
  HS65_GS_PAOI2X1 U655 ( .A(n1027), .B(n1026), .P(n1029), .Z(n1032) );
  HS65_GS_NAND2X2 U656 ( .A(n603), .B(n604), .Z(n601) );
  HS65_GS_OAI21X2 U657 ( .A(n603), .B(n604), .C(n601), .Z(n1033) );
  HS65_GS_NOR2X2 U658 ( .A(n1032), .B(n1033), .Z(n602) );
  HS65_GS_AOI12X2 U659 ( .A(n604), .B(n603), .C(n602), .Z(n1035) );
  HS65_GS_NAND2X2 U660 ( .A(n607), .B(n608), .Z(n605) );
  HS65_GS_OAI21X2 U661 ( .A(n607), .B(n608), .C(n605), .Z(n1036) );
  HS65_GS_NOR2X2 U662 ( .A(n1035), .B(n1036), .Z(n606) );
  HS65_GS_AOI12X2 U663 ( .A(n608), .B(n607), .C(n606), .Z(n1039) );
  HS65_GS_NAND2X2 U664 ( .A(n610), .B(n611), .Z(n609) );
  HS65_GS_OAI21X2 U665 ( .A(n610), .B(n611), .C(n609), .Z(n1038) );
  HS65_GS_NOR2X2 U666 ( .A(n1039), .B(n1038), .Z(n1037) );
  HS65_GS_AOI12X2 U667 ( .A(n611), .B(n610), .C(n1037), .Z(n1043) );
  HS65_GS_NAND2X2 U668 ( .A(n613), .B(n614), .Z(n612) );
  HS65_GS_OAI21X2 U669 ( .A(n613), .B(n614), .C(n612), .Z(n1042) );
  HS65_GS_NOR2X2 U670 ( .A(n1043), .B(n1042), .Z(n1041) );
  HS65_GS_AOI12X2 U671 ( .A(n614), .B(n613), .C(n1041), .Z(n1438) );
  HS65_GS_FA1X4 U672 ( .A0(\mul_a1/fa1_c1_r[26] ), .B0(n616), .CI(n615), .CO(
        n1441), .S0(n620) );
  HS65_GS_FA1X4 U673 ( .A0(\mul_a1/fa1_c1_r[25] ), .B0(n618), .CI(n617), .CO(
        n619), .S0(n613) );
  HS65_GS_NAND2X2 U674 ( .A(n620), .B(n619), .Z(n621) );
  HS65_GS_OAI21X2 U675 ( .A(n620), .B(n619), .C(n621), .Z(n1439) );
  HS65_GS_OAI21X2 U676 ( .A(n1438), .B(n1439), .C(n621), .Z(n1440) );
  HS65_GS_PAOI2X1 U677 ( .A(n1007), .B(n1006), .P(n1009), .Z(n1003) );
  HS65_GS_NOR2X2 U678 ( .A(n1004), .B(n1003), .Z(n622) );
  HS65_GSS_XOR3X2 U679 ( .A(n622), .B(\mul_a1/fa1_s1_r[33] ), .C(
        \mul_a1/fa1_c1_r[32] ), .Z(n623) );
  HS65_GSS_XOR3X2 U680 ( .A(n625), .B(n624), .C(n623), .Z(
        \mul_a1/result_sat[15] ) );
  HS65_GS_IVX2 U681 ( .A(y_z1[15]), .Z(n1483) );
  HS65_GS_IVX2 U682 ( .A(y_z1[14]), .Z(n1655) );
  HS65_GS_IVX2 U683 ( .A(y_z1[13]), .Z(n1657) );
  HS65_GS_IVX2 U684 ( .A(y_z1[12]), .Z(n1659) );
  HS65_GS_IVX2 U685 ( .A(y_z1[11]), .Z(n1661) );
  HS65_GS_IVX2 U686 ( .A(y_z1[10]), .Z(n1663) );
  HS65_GS_IVX2 U687 ( .A(y_z1[9]), .Z(n1665) );
  HS65_GS_IVX2 U688 ( .A(y_z1[8]), .Z(n1667) );
  HS65_GS_IVX2 U689 ( .A(y_z1[7]), .Z(n1669) );
  HS65_GS_IVX2 U690 ( .A(y_z1[6]), .Z(n1671) );
  HS65_GS_IVX2 U691 ( .A(y_z1[5]), .Z(n1673) );
  HS65_GS_IVX2 U692 ( .A(y_z1[4]), .Z(n1675) );
  HS65_GS_IVX2 U693 ( .A(y_z1[3]), .Z(n1677) );
  HS65_GS_IVX2 U694 ( .A(y_z1[2]), .Z(n1484) );
  HS65_GS_IVX2 U695 ( .A(y_z1[1]), .Z(n1447) );
  HS65_GS_IVX2 U696 ( .A(y_z1[0]), .Z(n1446) );
  HS65_GS_NOR2X2 U697 ( .A(y_z1[15]), .B(n1500), .Z(n1708) );
  HS65_GS_AND2X4 U698 ( .A(\mul_b0/fa1_s0_r[31] ), .B(\mul_b0/fa1_s1_r[31] ), 
        .Z(n627) );
  HS65_GSS_XOR2X3 U699 ( .A(\mul_b0/fa1_s0_r[32] ), .B(\mul_b0/fa1_s1_r[32] ), 
        .Z(n626) );
  HS65_GS_AND2X4 U700 ( .A(\mul_b0/fa1_s1_r[32] ), .B(\mul_b0/fa1_s0_r[32] ), 
        .Z(n742) );
  HS65_GS_AND2X4 U701 ( .A(\mul_b0/fa1_s0_r[29] ), .B(\mul_b0/fa1_s1_r[29] ), 
        .Z(n631) );
  HS65_GSS_XOR2X3 U702 ( .A(\mul_b0/fa1_s0_r[30] ), .B(\mul_b0/fa1_s1_r[30] ), 
        .Z(n630) );
  HS65_GSS_XOR2X3 U703 ( .A(\mul_b0/fa1_s0_r[31] ), .B(\mul_b0/fa1_s1_r[31] ), 
        .Z(n629) );
  HS65_GS_AND2X4 U704 ( .A(\mul_b0/fa1_s0_r[30] ), .B(\mul_b0/fa1_s1_r[30] ), 
        .Z(n628) );
  HS65_GS_FA1X4 U705 ( .A0(\mul_b0/fa1_s2_r[32] ), .B0(n627), .CI(n626), .CO(
        n743), .S0(n739) );
  HS65_GS_FA1X4 U706 ( .A0(\mul_b0/fa1_s2_r[31] ), .B0(n629), .CI(n628), .CO(
        n738), .S0(n735) );
  HS65_GSS_XNOR2X3 U707 ( .A(n739), .B(n738), .Z(n1054) );
  HS65_GS_IVX2 U708 ( .A(n1054), .Z(n737) );
  HS65_GS_AOI12X2 U709 ( .A(n734), .B(n735), .C(n737), .Z(n1053) );
  HS65_GS_NAND2X2 U710 ( .A(n735), .B(n734), .Z(n733) );
  HS65_GS_IVX2 U711 ( .A(n733), .Z(n736) );
  HS65_GS_AND2X4 U712 ( .A(\mul_b0/fa1_s0_r[28] ), .B(\mul_b0/fa1_s1_r[28] ), 
        .Z(n633) );
  HS65_GSS_XOR2X3 U713 ( .A(\mul_b0/fa1_s0_r[29] ), .B(\mul_b0/fa1_s1_r[29] ), 
        .Z(n632) );
  HS65_GS_FA1X4 U714 ( .A0(\mul_b0/fa1_s2_r[30] ), .B0(n631), .CI(n630), .CO(
        n734), .S0(n1061) );
  HS65_GS_AND2X4 U715 ( .A(\mul_b0/fa1_s0_r[27] ), .B(\mul_b0/fa1_s1_r[27] ), 
        .Z(n635) );
  HS65_GSS_XOR2X3 U716 ( .A(\mul_b0/fa1_s0_r[28] ), .B(\mul_b0/fa1_s1_r[28] ), 
        .Z(n634) );
  HS65_GS_FA1X4 U717 ( .A0(\mul_b0/fa1_s2_r[29] ), .B0(n633), .CI(n632), .CO(
        n1062), .S0(n1064) );
  HS65_GS_FA1X4 U718 ( .A0(\mul_b0/fa1_s2_r[28] ), .B0(n635), .CI(n634), .CO(
        n1065), .S0(n1508) );
  HS65_GSS_XOR2X3 U719 ( .A(\mul_b0/fa1_s0_r[27] ), .B(\mul_b0/fa1_s1_r[27] ), 
        .Z(n726) );
  HS65_GS_AND2X4 U720 ( .A(\mul_b0/fa1_s0_r[26] ), .B(\mul_b0/fa1_s1_r[26] ), 
        .Z(n725) );
  HS65_GS_AND2X4 U721 ( .A(\mul_b0/fa1_s0_r[24] ), .B(\mul_b0/fa1_s1_r[24] ), 
        .Z(n637) );
  HS65_GSS_XOR2X3 U722 ( .A(\mul_b0/fa1_s0_r[25] ), .B(\mul_b0/fa1_s1_r[25] ), 
        .Z(n636) );
  HS65_GS_AND2X4 U723 ( .A(\mul_b0/fa1_s1_r[25] ), .B(\mul_b0/fa1_s0_r[25] ), 
        .Z(n728) );
  HS65_GSS_XOR2X3 U724 ( .A(\mul_b0/fa1_s0_r[26] ), .B(\mul_b0/fa1_s1_r[26] ), 
        .Z(n727) );
  HS65_GSS_XOR2X3 U725 ( .A(\mul_b0/fa1_s0_r[24] ), .B(\mul_b0/fa1_s1_r[24] ), 
        .Z(n639) );
  HS65_GS_AND2X4 U726 ( .A(\mul_b0/fa1_s0_r[23] ), .B(\mul_b0/fa1_s1_r[23] ), 
        .Z(n638) );
  HS65_GS_FA1X4 U727 ( .A0(\mul_b0/fa1_s2_r[25] ), .B0(n637), .CI(n636), .CO(
        n724), .S0(n720) );
  HS65_GS_AND2X4 U728 ( .A(\mul_b0/fa1_s0_r[22] ), .B(\mul_b0/fa1_s1_r[22] ), 
        .Z(n641) );
  HS65_GSS_XOR2X3 U729 ( .A(\mul_b0/fa1_s0_r[23] ), .B(\mul_b0/fa1_s1_r[23] ), 
        .Z(n640) );
  HS65_GS_FA1X4 U730 ( .A0(\mul_b0/fa1_s2_r[24] ), .B0(n639), .CI(n638), .CO(
        n721), .S0(n717) );
  HS65_GSS_XOR2X3 U731 ( .A(\mul_b0/fa1_s0_r[22] ), .B(\mul_b0/fa1_s1_r[22] ), 
        .Z(n642) );
  HS65_GS_FA1X4 U732 ( .A0(\mul_b0/fa1_s2_r[23] ), .B0(n641), .CI(n640), .CO(
        n718), .S0(n714) );
  HS65_GS_FA1X4 U733 ( .A0(\mul_b0/fa1_s0_r[21] ), .B0(\mul_b0/fa1_s1_r[21] ), 
        .CI(\mul_b0/fa1_c0_r[20] ), .CO(n643), .S0(n644) );
  HS65_GS_FA1X4 U734 ( .A0(\mul_b0/fa1_s2_r[22] ), .B0(n643), .CI(n642), .CO(
        n715), .S0(n711) );
  HS65_GS_FA1X4 U735 ( .A0(\mul_b0/fa1_s0_r[20] ), .B0(\mul_b0/fa1_s1_r[20] ), 
        .CI(\mul_b0/fa1_c0_r[19] ), .CO(n645), .S0(n647) );
  HS65_GS_FA1X4 U736 ( .A0(\mul_b0/fa1_s2_r[21] ), .B0(n645), .CI(n644), .CO(
        n712), .S0(n708) );
  HS65_GS_FA1X4 U737 ( .A0(\mul_b0/fa1_s0_r[19] ), .B0(\mul_b0/fa1_s1_r[19] ), 
        .CI(\mul_b0/fa1_c0_r[18] ), .CO(n646), .S0(n648) );
  HS65_GS_FA1X4 U738 ( .A0(\mul_b0/fa1_s2_r[20] ), .B0(n647), .CI(n646), .CO(
        n709), .S0(n705) );
  HS65_GS_FA1X4 U739 ( .A0(\mul_b0/fa1_s0_r[18] ), .B0(\mul_b0/fa1_s1_r[18] ), 
        .CI(\mul_b0/fa1_c0_r[17] ), .CO(n649), .S0(n650) );
  HS65_GS_FA1X4 U740 ( .A0(\mul_b0/fa1_s2_r[19] ), .B0(n649), .CI(n648), .CO(
        n706), .S0(n702) );
  HS65_GS_FA1X4 U741 ( .A0(\mul_b0/fa1_s0_r[17] ), .B0(\mul_b0/fa1_s1_r[17] ), 
        .CI(\mul_b0/fa1_c0_r[16] ), .CO(n651), .S0(n652) );
  HS65_GS_FA1X4 U742 ( .A0(\mul_b0/fa1_s2_r[18] ), .B0(n651), .CI(n650), .CO(
        n703), .S0(n699) );
  HS65_GS_FA1X4 U743 ( .A0(\mul_b0/fa1_s0_r[16] ), .B0(\mul_b0/fa1_s1_r[16] ), 
        .CI(\mul_b0/fa1_c0_r[15] ), .CO(n653), .S0(n654) );
  HS65_GS_FA1X4 U744 ( .A0(\mul_b0/fa1_s2_r[17] ), .B0(n653), .CI(n652), .CO(
        n700), .S0(n695) );
  HS65_GS_FA1X4 U745 ( .A0(\mul_b0/fa1_s0_r[15] ), .B0(\mul_b0/fa1_s1_r[15] ), 
        .CI(\mul_b0/fa1_c0_r[14] ), .CO(n655), .S0(n657) );
  HS65_GS_FA1X4 U746 ( .A0(\mul_b0/fa1_s2_r[16] ), .B0(n655), .CI(n654), .CO(
        n696), .S0(n692) );
  HS65_GS_NAND2X2 U747 ( .A(n692), .B(n693), .Z(n656) );
  HS65_GS_OAI21X2 U748 ( .A(n692), .B(n693), .C(n656), .Z(n1081) );
  HS65_GS_FA1X4 U749 ( .A0(\mul_b0/fa1_s0_r[14] ), .B0(\mul_b0/fa1_s1_r[14] ), 
        .CI(\mul_b0/fa1_c0_r[13] ), .CO(n658), .S0(n660) );
  HS65_GS_FA1X4 U750 ( .A0(\mul_b0/fa1_s2_r[15] ), .B0(n658), .CI(n657), .CO(
        n693), .S0(n690) );
  HS65_GS_NOR2X2 U751 ( .A(n691), .B(n690), .Z(n659) );
  HS65_GS_AOI12X2 U752 ( .A(n690), .B(n691), .C(n659), .Z(n1078) );
  HS65_GS_FA1X4 U753 ( .A0(\mul_b0/fa1_s0_r[13] ), .B0(\mul_b0/fa1_s1_r[13] ), 
        .CI(\mul_b0/fa1_c0_r[12] ), .CO(n661), .S0(n662) );
  HS65_GS_FA1X4 U754 ( .A0(\mul_b0/fa1_s2_r[14] ), .B0(n661), .CI(n660), .CO(
        n691), .S0(n687) );
  HS65_GS_FA1X4 U755 ( .A0(\mul_b0/fa1_s2_r[13] ), .B0(n663), .CI(n662), .CO(
        n688), .S0(n685) );
  HS65_GS_FA1X4 U756 ( .A0(\mul_b0/fa1_s0_r[12] ), .B0(\mul_b0/fa1_s1_r[12] ), 
        .CI(\mul_b0/fa1_c0_r[11] ), .CO(n663), .S0(n677) );
  HS65_GS_FA1X4 U757 ( .A0(\mul_b0/fa1_s0_r[11] ), .B0(\mul_b0/fa1_s1_r[11] ), 
        .CI(\mul_b0/fa1_c0_r[10] ), .CO(n678), .S0(n682) );
  HS65_GS_FA1X4 U758 ( .A0(\mul_b0/fa1_s0_r[10] ), .B0(\mul_b0/fa1_s1_r[10] ), 
        .CI(\mul_b0/fa1_c0_r[9] ), .CO(n681), .S0(n675) );
  HS65_GS_OR2X4 U759 ( .A(n681), .B(n682), .Z(n674) );
  HS65_GS_OAI22X1 U760 ( .A(n681), .B(n682), .C(n676), .D(n675), .Z(n672) );
  HS65_GS_FA1X4 U761 ( .A0(\mul_b0/fa1_s0_r[9] ), .B0(\mul_b0/fa1_s1_r[9] ), 
        .CI(\mul_b0/fa1_c0_r[8] ), .CO(n676), .S0(n670) );
  HS65_GS_NOR2X2 U762 ( .A(\mul_b0/fa1_c0_r[6] ), .B(\mul_b0/fa1_s0_r[7] ), 
        .Z(n665) );
  HS65_GS_NAND2X2 U763 ( .A(\mul_b0/fa1_c0_r[5] ), .B(\mul_b0/fa1_s0_r[6] ), 
        .Z(n664) );
  HS65_GS_NOR2X2 U764 ( .A(n665), .B(n664), .Z(n667) );
  HS65_GS_CB4I1X4 U765 ( .A(\mul_b0/fa1_c0_r[6] ), .B(\mul_b0/fa1_s0_r[7] ), 
        .C(n667), .D(n666), .Z(n669) );
  HS65_GS_FA1X4 U766 ( .A0(\mul_b0/fa1_s0_r[8] ), .B0(\mul_b0/fa1_s1_r[8] ), 
        .CI(\mul_b0/fa1_c0_r[7] ), .CO(n668), .S0(n666) );
  HS65_GS_PAOI2X1 U767 ( .A(n670), .B(n669), .P(n668), .Z(n671) );
  HS65_GS_NOR2X2 U768 ( .A(n672), .B(n671), .Z(n673) );
  HS65_GS_AO31X4 U769 ( .A(n676), .B(n675), .C(n674), .D(n673), .Z(n680) );
  HS65_GS_FA1X4 U770 ( .A0(\mul_b0/fa1_s2_r[12] ), .B0(n678), .CI(n677), .CO(
        n684), .S0(n679) );
  HS65_GS_CB4I1X4 U771 ( .A(n682), .B(n681), .C(n680), .D(n679), .Z(n683) );
  HS65_GS_PAOI2X1 U772 ( .A(n685), .B(n684), .P(n683), .Z(n1074) );
  HS65_GS_NAND2X2 U773 ( .A(n687), .B(n688), .Z(n686) );
  HS65_GS_OAI21X2 U774 ( .A(n687), .B(n688), .C(n686), .Z(n1073) );
  HS65_GS_NOR2X2 U775 ( .A(n1074), .B(n1073), .Z(n1072) );
  HS65_GS_AOI12X2 U776 ( .A(n688), .B(n687), .C(n1072), .Z(n1077) );
  HS65_GS_NAND2X2 U777 ( .A(n1078), .B(n1077), .Z(n689) );
  HS65_GS_OAI21X2 U778 ( .A(n691), .B(n690), .C(n689), .Z(n1080) );
  HS65_GS_NOR2X2 U779 ( .A(n1081), .B(n1080), .Z(n1079) );
  HS65_GS_AOI12X2 U780 ( .A(n693), .B(n692), .C(n1079), .Z(n1085) );
  HS65_GS_NAND2X2 U781 ( .A(n695), .B(n696), .Z(n694) );
  HS65_GS_OAI21X2 U782 ( .A(n695), .B(n696), .C(n694), .Z(n1084) );
  HS65_GS_NOR2X2 U783 ( .A(n1085), .B(n1084), .Z(n1083) );
  HS65_GS_AOI12X2 U784 ( .A(n696), .B(n695), .C(n1083), .Z(n1089) );
  HS65_GS_NOR2X2 U785 ( .A(n700), .B(n699), .Z(n697) );
  HS65_GS_AOI12X2 U786 ( .A(n699), .B(n700), .C(n697), .Z(n1088) );
  HS65_GS_NAND2X2 U787 ( .A(n1089), .B(n1088), .Z(n698) );
  HS65_GS_OAI21X2 U788 ( .A(n700), .B(n699), .C(n698), .Z(n1092) );
  HS65_GS_NAND2X2 U789 ( .A(n702), .B(n703), .Z(n701) );
  HS65_GS_OAI21X2 U790 ( .A(n702), .B(n703), .C(n701), .Z(n1091) );
  HS65_GS_NOR2X2 U791 ( .A(n1092), .B(n1091), .Z(n1090) );
  HS65_GS_AOI12X2 U792 ( .A(n703), .B(n702), .C(n1090), .Z(n1096) );
  HS65_GS_NAND2X2 U793 ( .A(n705), .B(n706), .Z(n704) );
  HS65_GS_OAI21X2 U794 ( .A(n705), .B(n706), .C(n704), .Z(n1095) );
  HS65_GS_NOR2X2 U795 ( .A(n1096), .B(n1095), .Z(n1094) );
  HS65_GS_AOI12X2 U796 ( .A(n706), .B(n705), .C(n1094), .Z(n1100) );
  HS65_GS_NAND2X2 U797 ( .A(n708), .B(n709), .Z(n707) );
  HS65_GS_OAI21X2 U798 ( .A(n708), .B(n709), .C(n707), .Z(n1099) );
  HS65_GS_NOR2X2 U799 ( .A(n1100), .B(n1099), .Z(n1098) );
  HS65_GS_AOI12X2 U800 ( .A(n709), .B(n708), .C(n1098), .Z(n1104) );
  HS65_GS_NAND2X2 U801 ( .A(n711), .B(n712), .Z(n710) );
  HS65_GS_OAI21X2 U802 ( .A(n711), .B(n712), .C(n710), .Z(n1103) );
  HS65_GS_NOR2X2 U803 ( .A(n1104), .B(n1103), .Z(n1102) );
  HS65_GS_AOI12X2 U804 ( .A(n712), .B(n711), .C(n1102), .Z(n1108) );
  HS65_GS_NAND2X2 U805 ( .A(n714), .B(n715), .Z(n713) );
  HS65_GS_OAI21X2 U806 ( .A(n714), .B(n715), .C(n713), .Z(n1107) );
  HS65_GS_NOR2X2 U807 ( .A(n1108), .B(n1107), .Z(n1106) );
  HS65_GS_AOI12X2 U808 ( .A(n715), .B(n714), .C(n1106), .Z(n1112) );
  HS65_GS_NAND2X2 U809 ( .A(n717), .B(n718), .Z(n716) );
  HS65_GS_OAI21X2 U810 ( .A(n717), .B(n718), .C(n716), .Z(n1111) );
  HS65_GS_NOR2X2 U811 ( .A(n1112), .B(n1111), .Z(n1110) );
  HS65_GS_AOI12X2 U812 ( .A(n718), .B(n717), .C(n1110), .Z(n1116) );
  HS65_GS_NAND2X2 U813 ( .A(n720), .B(n721), .Z(n719) );
  HS65_GS_OAI21X2 U814 ( .A(n720), .B(n721), .C(n719), .Z(n1115) );
  HS65_GS_NOR2X2 U815 ( .A(n1116), .B(n1115), .Z(n1114) );
  HS65_GS_AOI12X2 U816 ( .A(n721), .B(n720), .C(n1114), .Z(n1120) );
  HS65_GS_NAND2X2 U817 ( .A(n723), .B(n724), .Z(n722) );
  HS65_GS_OAI21X2 U818 ( .A(n723), .B(n724), .C(n722), .Z(n1119) );
  HS65_GS_NOR2X2 U819 ( .A(n1120), .B(n1119), .Z(n1118) );
  HS65_GS_AOI12X2 U820 ( .A(n724), .B(n723), .C(n1118), .Z(n1504) );
  HS65_GS_FA1X4 U821 ( .A0(\mul_b0/fa1_s2_r[27] ), .B0(n726), .CI(n725), .CO(
        n1507), .S0(n730) );
  HS65_GS_FA1X4 U822 ( .A0(\mul_b0/fa1_s2_r[26] ), .B0(n728), .CI(n727), .CO(
        n729), .S0(n723) );
  HS65_GS_NAND2X2 U823 ( .A(n730), .B(n729), .Z(n731) );
  HS65_GS_OAI21X2 U824 ( .A(n730), .B(n729), .C(n731), .Z(n1505) );
  HS65_GS_OAI21X2 U825 ( .A(n1504), .B(n1505), .C(n731), .Z(n1506) );
  HS65_GS_IVX2 U826 ( .A(n732), .Z(n1059) );
  HS65_GS_OAI21X2 U827 ( .A(n735), .B(n734), .C(n733), .Z(n1058) );
  HS65_GS_NOR2X2 U828 ( .A(n1059), .B(n1058), .Z(n1057) );
  HS65_GS_AOI12X2 U829 ( .A(n737), .B(n736), .C(n1057), .Z(n1056) );
  HS65_GS_NAND2X2 U830 ( .A(n739), .B(n738), .Z(n740) );
  HS65_GS_OAI21X2 U831 ( .A(n1053), .B(n1056), .C(n740), .Z(n741) );
  HS65_GSS_XOR3X2 U832 ( .A(n743), .B(n742), .C(n741), .Z(n744) );
  HS65_GSS_XOR2X3 U833 ( .A(\mul_b0/fa1_s2_r[33] ), .B(n744), .Z(n745) );
  HS65_GSS_XOR3X2 U834 ( .A(\mul_b0/fa1_s0_r[33] ), .B(\mul_b0/fa1_s1_r[33] ), 
        .C(n745), .Z(\mul_b0/result_sat[15] ) );
  HS65_GS_IVX2 U835 ( .A(x_z1[15]), .Z(n1554) );
  HS65_GS_AND2X4 U836 ( .A(p_b1[1]), .B(p_b0[1]), .Z(n785) );
  HS65_GSS_XOR2X3 U837 ( .A(p_b1[1]), .B(p_b0[1]), .Z(n788) );
  HS65_GS_FA1X4 U838 ( .A0(p_b0[2]), .B0(p_b1[2]), .CI(p_b2[2]), .CO(n781), 
        .S0(n783) );
  HS65_GS_FA1X4 U839 ( .A0(p_b0[3]), .B0(p_b1[3]), .CI(p_b2[3]), .CO(n777), 
        .S0(n779) );
  HS65_GS_FA1X4 U840 ( .A0(p_b0[4]), .B0(p_b1[4]), .CI(p_b2[4]), .CO(n773), 
        .S0(n775) );
  HS65_GS_FA1X4 U841 ( .A0(p_b0[5]), .B0(p_b1[5]), .CI(p_b2[5]), .CO(n769), 
        .S0(n771) );
  HS65_GS_FA1X4 U842 ( .A0(p_b0[6]), .B0(p_b1[6]), .CI(p_b2[6]), .CO(n765), 
        .S0(n767) );
  HS65_GS_FA1X4 U843 ( .A0(p_b0[7]), .B0(p_b1[7]), .CI(p_b2[7]), .CO(n761), 
        .S0(n763) );
  HS65_GS_FA1X4 U844 ( .A0(p_b0[8]), .B0(p_b1[8]), .CI(p_b2[8]), .CO(n753), 
        .S0(n759) );
  HS65_GS_FA1X4 U845 ( .A0(p_b0[9]), .B0(p_b1[9]), .CI(p_b2[9]), .CO(n757), 
        .S0(n751) );
  HS65_GS_FA1X4 U846 ( .A0(p_b0[10]), .B0(p_b1[10]), .CI(p_b2[10]), .CO(n749), 
        .S0(n755) );
  HS65_GS_FA1X4 U847 ( .A0(p_b0[11]), .B0(p_b1[11]), .CI(p_b2[11]), .CO(n831), 
        .S0(n747) );
  HS65_GS_IVX2 U848 ( .A(n746), .Z(n828) );
  HS65_GS_FA1X4 U849 ( .A0(n749), .B0(n748), .CI(n747), .CO(n830), .S0(n750)
         );
  HS65_GS_IVX2 U850 ( .A(n750), .Z(n827) );
  HS65_GS_FA1X4 U851 ( .A0(n753), .B0(n752), .CI(n751), .CO(n756), .S0(n754)
         );
  HS65_GS_IVX2 U852 ( .A(n754), .Z(n820) );
  HS65_GS_FA1X4 U853 ( .A0(n757), .B0(n756), .CI(n755), .CO(n748), .S0(n758)
         );
  HS65_GS_IVX2 U854 ( .A(n758), .Z(n824) );
  HS65_GS_FA1X4 U855 ( .A0(n761), .B0(n760), .CI(n759), .CO(n752), .S0(n762)
         );
  HS65_GS_IVX2 U856 ( .A(n762), .Z(n816) );
  HS65_GS_FA1X4 U857 ( .A0(n765), .B0(n764), .CI(n763), .CO(n760), .S0(n766)
         );
  HS65_GS_IVX2 U858 ( .A(n766), .Z(n812) );
  HS65_GS_FA1X4 U859 ( .A0(n769), .B0(n768), .CI(n767), .CO(n764), .S0(n770)
         );
  HS65_GS_IVX2 U860 ( .A(n770), .Z(n808) );
  HS65_GS_FA1X4 U861 ( .A0(n773), .B0(n772), .CI(n771), .CO(n768), .S0(n774)
         );
  HS65_GS_IVX2 U862 ( .A(n774), .Z(n804) );
  HS65_GS_FA1X4 U863 ( .A0(n777), .B0(n776), .CI(n775), .CO(n772), .S0(n778)
         );
  HS65_GS_IVX2 U864 ( .A(n778), .Z(n800) );
  HS65_GS_FA1X4 U865 ( .A0(n781), .B0(n780), .CI(n779), .CO(n776), .S0(n782)
         );
  HS65_GS_IVX2 U866 ( .A(n782), .Z(n796) );
  HS65_GS_FA1X4 U867 ( .A0(n785), .B0(n784), .CI(n783), .CO(n780), .S0(n786)
         );
  HS65_GS_IVX2 U868 ( .A(n786), .Z(n791) );
  HS65_GS_FA1X4 U869 ( .A0(p_b2[1]), .B0(n788), .CI(n787), .CO(n784), .S0(n789) );
  HS65_GS_IVX2 U870 ( .A(n789), .Z(n793) );
  HS65_GS_FA1X4 U871 ( .A0(p_b2[0]), .B0(p_b0[0]), .CI(p_b1[0]), .CO(n787), 
        .S0(n790) );
  HS65_GS_IVX2 U872 ( .A(n790), .Z(n922) );
  HS65_GS_NAND2X2 U873 ( .A(n1249), .B(p_a1[1]), .Z(n1248) );
  HS65_GS_NAND3AX3 U874 ( .A(n1248), .B(p_a2[1]), .C(n793), .Z(n795) );
  HS65_GS_FA1X4 U875 ( .A0(p_a2[2]), .B0(p_a1[2]), .CI(n791), .CO(n798), .S0(
        n1253) );
  HS65_GS_FA1X4 U876 ( .A0(p_a2[1]), .B0(n793), .CI(n792), .CO(n794), .S0(
        n1249) );
  HS65_GS_CB4I1X4 U877 ( .A(p_a1[1]), .B(n1249), .C(n794), .D(n795), .Z(n1252)
         );
  HS65_GS_NAND2X2 U878 ( .A(n1253), .B(n1252), .Z(n1251) );
  HS65_GS_NAND2X2 U879 ( .A(n795), .B(n1251), .Z(n797) );
  HS65_GS_NOR2X2 U880 ( .A(n798), .B(n797), .Z(n799) );
  HS65_GS_FA1X4 U881 ( .A0(p_a2[3]), .B0(p_a1[3]), .CI(n796), .CO(n802), .S0(
        n1257) );
  HS65_GSS_XNOR2X3 U882 ( .A(n798), .B(n797), .Z(n1256) );
  HS65_GS_NOR2X2 U883 ( .A(n1257), .B(n1256), .Z(n1255) );
  HS65_GS_NOR2X2 U884 ( .A(n799), .B(n1255), .Z(n801) );
  HS65_GS_NAND2X2 U885 ( .A(n802), .B(n801), .Z(n803) );
  HS65_GS_FA1X4 U886 ( .A0(p_a2[4]), .B0(p_a1[4]), .CI(n800), .CO(n805), .S0(
        n1261) );
  HS65_GSS_XOR2X3 U887 ( .A(n802), .B(n801), .Z(n1260) );
  HS65_GS_NAND2X2 U888 ( .A(n1261), .B(n1260), .Z(n1259) );
  HS65_GS_NAND2X2 U889 ( .A(n803), .B(n1259), .Z(n806) );
  HS65_GS_NAND2X2 U890 ( .A(n805), .B(n806), .Z(n807) );
  HS65_GS_FA1X4 U891 ( .A0(p_a2[5]), .B0(p_a1[5]), .CI(n804), .CO(n809), .S0(
        n1265) );
  HS65_GSS_XOR2X3 U892 ( .A(n806), .B(n805), .Z(n1264) );
  HS65_GS_NAND2X2 U893 ( .A(n1265), .B(n1264), .Z(n1263) );
  HS65_GS_NAND2X2 U894 ( .A(n807), .B(n1263), .Z(n810) );
  HS65_GS_NAND2X2 U895 ( .A(n809), .B(n810), .Z(n811) );
  HS65_GS_FA1X4 U896 ( .A0(p_a2[6]), .B0(p_a1[6]), .CI(n808), .CO(n813), .S0(
        n1269) );
  HS65_GSS_XOR2X3 U897 ( .A(n810), .B(n809), .Z(n1268) );
  HS65_GS_NAND2X2 U898 ( .A(n1269), .B(n1268), .Z(n1267) );
  HS65_GS_NAND2X2 U899 ( .A(n811), .B(n1267), .Z(n814) );
  HS65_GS_NAND2X2 U900 ( .A(n813), .B(n814), .Z(n815) );
  HS65_GS_FA1X4 U901 ( .A0(p_a2[7]), .B0(p_a1[7]), .CI(n812), .CO(n817), .S0(
        n1273) );
  HS65_GSS_XOR2X3 U902 ( .A(n814), .B(n813), .Z(n1272) );
  HS65_GS_NAND2X2 U903 ( .A(n1273), .B(n1272), .Z(n1271) );
  HS65_GS_NAND2X2 U904 ( .A(n815), .B(n1271), .Z(n818) );
  HS65_GS_NAND2X2 U905 ( .A(n817), .B(n818), .Z(n819) );
  HS65_GS_FA1X4 U906 ( .A0(p_a2[8]), .B0(p_a1[8]), .CI(n816), .CO(n821), .S0(
        n1277) );
  HS65_GSS_XOR2X3 U907 ( .A(n818), .B(n817), .Z(n1276) );
  HS65_GS_NAND2X2 U908 ( .A(n1277), .B(n1276), .Z(n1275) );
  HS65_GS_NAND2X2 U909 ( .A(n819), .B(n1275), .Z(n822) );
  HS65_GS_NAND2X2 U910 ( .A(n821), .B(n822), .Z(n823) );
  HS65_GS_FA1X4 U911 ( .A0(p_a2[9]), .B0(p_a1[9]), .CI(n820), .CO(n1283), .S0(
        n1281) );
  HS65_GSS_XOR2X3 U912 ( .A(n822), .B(n821), .Z(n1280) );
  HS65_GS_NAND2X2 U913 ( .A(n1281), .B(n1280), .Z(n1279) );
  HS65_GS_NAND2X2 U914 ( .A(n823), .B(n1279), .Z(n1284) );
  HS65_GS_PAO2X4 U915 ( .A(n1283), .B(n1286), .P(n1284), .Z(n825) );
  HS65_GS_FA1X4 U916 ( .A0(p_a2[10]), .B0(p_a1[10]), .CI(n824), .CO(n826), 
        .S0(n1286) );
  HS65_GSS_XOR2X3 U917 ( .A(n825), .B(n826), .Z(n1295) );
  HS65_GS_AO22X4 U918 ( .A(n1294), .B(n1295), .C(n826), .D(n825), .Z(n1300) );
  HS65_GS_FA1X4 U919 ( .A0(p_a2[11]), .B0(p_a1[11]), .CI(n827), .CO(n1299), 
        .S0(n1294) );
  HS65_GS_FA1X4 U920 ( .A0(p_a2[12]), .B0(p_a1[12]), .CI(n828), .CO(n927), 
        .S0(n1298) );
  HS65_GS_FA1X4 U921 ( .A0(p_b0[12]), .B0(p_b1[12]), .CI(p_b2[12]), .CO(n836), 
        .S0(n829) );
  HS65_GS_FA1X4 U922 ( .A0(n831), .B0(n830), .CI(n829), .CO(n835), .S0(n746)
         );
  HS65_GS_IVX2 U923 ( .A(n832), .Z(n833) );
  HS65_GS_FA1X4 U924 ( .A0(p_a1[13]), .B0(p_a2[13]), .CI(n833), .CO(n843), 
        .S0(n925) );
  HS65_GS_FA1X4 U925 ( .A0(p_b0[13]), .B0(p_b1[13]), .CI(p_b2[13]), .CO(n840), 
        .S0(n834) );
  HS65_GS_FA1X4 U926 ( .A0(n836), .B0(n835), .CI(n834), .CO(n839), .S0(n832)
         );
  HS65_GS_IVX2 U927 ( .A(n837), .Z(n845) );
  HS65_GS_FA1X4 U928 ( .A0(p_b0[14]), .B0(p_b1[14]), .CI(p_b2[14]), .CO(n850), 
        .S0(n838) );
  HS65_GS_FA1X4 U929 ( .A0(n840), .B0(n839), .CI(n838), .CO(n849), .S0(n837)
         );
  HS65_GS_IVX2 U930 ( .A(p_b0[15]), .Z(n851) );
  HS65_GS_NAND2X2 U931 ( .A(p_b2[15]), .B(p_b1[15]), .Z(n852) );
  HS65_GS_OAI21X2 U932 ( .A(p_b2[15]), .B(p_b1[15]), .C(n852), .Z(n841) );
  HS65_GS_MUXI21X2 U933 ( .D0(p_b0[15]), .D1(n851), .S0(n841), .Z(n848) );
  HS65_GS_FA1X4 U934 ( .A0(n844), .B0(n843), .CI(n842), .CO(n857), .S0(n870)
         );
  HS65_GS_FA1X4 U935 ( .A0(p_a1[14]), .B0(p_a2[14]), .CI(n845), .CO(n856), 
        .S0(n842) );
  HS65_GS_FA1X4 U936 ( .A0(p_a1[15]), .B0(p_a2[15]), .CI(n846), .CO(n861), 
        .S0(n847) );
  HS65_GS_IVX2 U937 ( .A(n847), .Z(n855) );
  HS65_GS_FA1X4 U938 ( .A0(n850), .B0(n849), .CI(n848), .CO(n854), .S0(n846)
         );
  HS65_GS_OAI32X2 U939 ( .A(p_b0[15]), .B(p_b2[15]), .C(p_b1[15]), .D(n852), 
        .E(n851), .Z(n853) );
  HS65_GSS_XNOR2X3 U940 ( .A(n854), .B(n853), .Z(n858) );
  HS65_GSS_XNOR2X3 U941 ( .A(n859), .B(n858), .Z(n860) );
  HS65_GS_NAND2X2 U942 ( .A(n861), .B(n860), .Z(n863) );
  HS65_GS_FA1X4 U943 ( .A0(n857), .B0(n856), .CI(n855), .CO(n859), .S0(n868)
         );
  HS65_GS_NAND2X2 U944 ( .A(n859), .B(n858), .Z(n862) );
  HS65_GS_IVX2 U945 ( .A(valid_T3), .Z(n1706) );
  HS65_GS_NOR2X2 U946 ( .A(n861), .B(n860), .Z(n865) );
  HS65_GS_NOR3AX2 U947 ( .A(n862), .B(n1706), .C(n865), .Z(n1704) );
  HS65_GS_IVX2 U948 ( .A(n1704), .Z(n866) );
  HS65_GS_AOI12X2 U949 ( .A(n863), .B(n868), .C(n866), .Z(n1301) );
  HS65_GS_IVX2 U950 ( .A(n1301), .Z(n1291) );
  HS65_GS_IVX2 U951 ( .A(n863), .Z(n864) );
  HS65_GS_OAI21X2 U952 ( .A(n865), .B(n864), .C(valid_T3), .Z(n867) );
  HS65_GS_OAI12X3 U953 ( .A(n868), .B(n867), .C(n866), .Z(n1292) );
  HS65_GS_IVX2 U954 ( .A(n1292), .Z(n1304) );
  HS65_GS_NAND2X2 U955 ( .A(data_out[14]), .B(n1706), .Z(n869) );
  HS65_GS_CBI4I1X3 U956 ( .A(n870), .B(n1291), .C(n1304), .D(n869), .Z(n1766)
         );
  HS65_GS_IVX2 U957 ( .A(y_z2[14]), .Z(n1343) );
  HS65_GS_IVX2 U958 ( .A(y_z2[13]), .Z(n1341) );
  HS65_GS_IVX2 U959 ( .A(y_z2[12]), .Z(n1339) );
  HS65_GS_IVX2 U960 ( .A(y_z2[11]), .Z(n1337) );
  HS65_GS_IVX2 U961 ( .A(y_z2[10]), .Z(n1335) );
  HS65_GS_IVX2 U962 ( .A(y_z2[9]), .Z(n1333) );
  HS65_GS_IVX2 U963 ( .A(y_z2[8]), .Z(n1331) );
  HS65_GS_IVX2 U964 ( .A(y_z2[7]), .Z(n1329) );
  HS65_GS_IVX2 U965 ( .A(y_z2[6]), .Z(n1327) );
  HS65_GS_IVX2 U966 ( .A(y_z2[5]), .Z(n1325) );
  HS65_GS_IVX2 U967 ( .A(y_z2[4]), .Z(n1323) );
  HS65_GS_IVX2 U968 ( .A(y_z2[3]), .Z(n1321) );
  HS65_GS_IVX2 U969 ( .A(y_z2[2]), .Z(n1319) );
  HS65_GS_IVX2 U970 ( .A(y_z2[1]), .Z(n1317) );
  HS65_GS_IVX2 U971 ( .A(y_z2[0]), .Z(n1247) );
  HS65_GS_NOR2X2 U972 ( .A(y_z2[15]), .B(n1182), .Z(n1707) );
  HS65_GS_IVX2 U973 ( .A(y_z2[15]), .Z(n1346) );
  HS65_GS_HA1X4 U974 ( .A0(n1346), .B0(n871), .S0(n872) );
  HS65_GSS_XOR2X3 U975 ( .A(n1707), .B(n872), .Z(\mul_a2/fa1_s1[25] ) );
  HS65_GS_MUXI21X2 U976 ( .D0(n874), .D1(n873), .S0(n1191), .Z(n895) );
  HS65_GS_FA1X4 U977 ( .A0(n877), .B0(n876), .CI(n875), .CO(n885), .S0(n892)
         );
  HS65_GS_FA1X4 U978 ( .A0(n880), .B0(n879), .CI(n878), .CO(n876), .S0(n890)
         );
  HS65_GS_FA1X4 U979 ( .A0(n883), .B0(n882), .CI(n881), .CO(n415), .S0(n889)
         );
  HS65_GS_FA1X4 U980 ( .A0(n886), .B0(n885), .CI(n884), .CO(n882), .S0(n888)
         );
  HS65_GS_OR3X4 U981 ( .A(n890), .B(n889), .C(n888), .Z(n887) );
  HS65_GS_OAI21X2 U982 ( .A(n892), .B(n887), .C(\mul_a2/result_sat[15] ), .Z(
        n1216) );
  HS65_GS_OAI21X2 U983 ( .A(n894), .B(n895), .C(n1216), .Z(n893) );
  HS65_GS_AND3X4 U984 ( .A(n890), .B(n889), .C(n888), .Z(n891) );
  HS65_GS_AOI12X2 U985 ( .A(n892), .B(n891), .C(\mul_a2/result_sat[15] ), .Z(
        n1215) );
  HS65_GS_IVX2 U986 ( .A(n1215), .Z(n1702) );
  HS65_GS_CBI4I1X3 U987 ( .A(n895), .B(n894), .C(n893), .D(n1702), .Z(
        \mul_a2/result_sat[2] ) );
  HS65_GSS_XNOR2X3 U988 ( .A(n897), .B(n896), .Z(n900) );
  HS65_GS_OAI21X2 U989 ( .A(n899), .B(n900), .C(n1216), .Z(n898) );
  HS65_GS_CBI4I1X3 U990 ( .A(n900), .B(n899), .C(n898), .D(n1702), .Z(
        \mul_a2/result_sat[5] ) );
  HS65_GSS_XNOR2X3 U991 ( .A(n902), .B(n901), .Z(n905) );
  HS65_GS_OAI21X2 U992 ( .A(n904), .B(n905), .C(n1216), .Z(n903) );
  HS65_GS_CBI4I1X3 U993 ( .A(n905), .B(n904), .C(n903), .D(n1702), .Z(
        \mul_a2/result_sat[7] ) );
  HS65_GSS_XNOR2X3 U994 ( .A(n907), .B(n906), .Z(n910) );
  HS65_GS_OAI21X2 U995 ( .A(n909), .B(n910), .C(n1216), .Z(n908) );
  HS65_GS_CBI4I1X3 U996 ( .A(n910), .B(n909), .C(n908), .D(n1702), .Z(
        \mul_a2/result_sat[8] ) );
  HS65_GSS_XNOR2X3 U997 ( .A(n912), .B(n911), .Z(n915) );
  HS65_GS_OAI21X2 U998 ( .A(n914), .B(n915), .C(n1216), .Z(n913) );
  HS65_GS_CBI4I1X3 U999 ( .A(n915), .B(n914), .C(n913), .D(n1702), .Z(
        \mul_a2/result_sat[9] ) );
  HS65_GSS_XNOR2X3 U1000 ( .A(n917), .B(n916), .Z(n921) );
  HS65_GS_IVX2 U1001 ( .A(n918), .Z(n920) );
  HS65_GS_OAI21X2 U1002 ( .A(n920), .B(n921), .C(n1216), .Z(n919) );
  HS65_GS_CBI4I1X3 U1003 ( .A(n921), .B(n920), .C(n919), .D(n1702), .Z(
        \mul_a2/result_sat[12] ) );
  HS65_GS_MUX21I1X3 U1004 ( .D0(n1446), .D1(data_out[0]), .S0(n1305), .Z(n1809) );
  HS65_GS_FA1X4 U1005 ( .A0(p_a2[0]), .B0(p_a1[0]), .CI(n922), .CO(n792), .S0(
        n924) );
  HS65_GS_NAND2X2 U1006 ( .A(data_out[0]), .B(n1706), .Z(n923) );
  HS65_GS_CBI4I1X3 U1007 ( .A(n924), .B(n1291), .C(n1304), .D(n923), .Z(n1808)
         );
  HS65_GS_MUX21I1X3 U1008 ( .D0(n1447), .D1(data_out[1]), .S0(n1714), .Z(n1806) );
  HS65_GS_MUX21I1X3 U1009 ( .D0(n1484), .D1(data_out[2]), .S0(valid_in), .Z(
        n1803) );
  HS65_GS_MUX21I1X3 U1010 ( .D0(n1677), .D1(data_out[3]), .S0(valid_in), .Z(
        n1800) );
  HS65_GS_MUX21I1X3 U1011 ( .D0(n1675), .D1(data_out[4]), .S0(valid_in), .Z(
        n1797) );
  HS65_GS_MUX21I1X3 U1012 ( .D0(n1673), .D1(data_out[5]), .S0(valid_in), .Z(
        n1794) );
  HS65_GS_MUX21I1X3 U1013 ( .D0(n1671), .D1(data_out[6]), .S0(valid_in), .Z(
        n1791) );
  HS65_GS_MUX21I1X3 U1014 ( .D0(n1669), .D1(data_out[7]), .S0(valid_in), .Z(
        n1788) );
  HS65_GS_MUX21I1X3 U1015 ( .D0(n1667), .D1(data_out[8]), .S0(valid_in), .Z(
        n1785) );
  HS65_GS_MUX21I1X3 U1016 ( .D0(n1665), .D1(data_out[9]), .S0(valid_in), .Z(
        n1782) );
  HS65_GS_BFX4 U1017 ( .A(n1714), .Z(n1290) );
  HS65_GS_MUX21I1X3 U1018 ( .D0(n1659), .D1(data_out[12]), .S0(n1290), .Z(
        n1773) );
  HS65_GS_MUX21I1X3 U1019 ( .D0(n1657), .D1(data_out[13]), .S0(n1290), .Z(
        n1770) );
  HS65_GS_FA1X4 U1020 ( .A0(n927), .B0(n926), .CI(n925), .CO(n844), .S0(n929)
         );
  HS65_GS_NAND2X2 U1021 ( .A(data_out[13]), .B(n1706), .Z(n928) );
  HS65_GS_CBI4I1X3 U1022 ( .A(n929), .B(n1291), .C(n1304), .D(n928), .Z(n1769)
         );
  HS65_GS_MUX21I1X3 U1023 ( .D0(n1655), .D1(data_out[14]), .S0(n1290), .Z(
        n1767) );
  HS65_GS_IVX2 U1024 ( .A(x_z2[15]), .Z(n1693) );
  HS65_GS_IVX2 U1025 ( .A(x_z2[14]), .Z(n1692) );
  HS65_GS_IVX2 U1026 ( .A(x_z2[13]), .Z(n1691) );
  HS65_GS_IVX2 U1027 ( .A(x_z2[12]), .Z(n1690) );
  HS65_GS_IVX2 U1028 ( .A(x_z2[11]), .Z(n1689) );
  HS65_GS_IVX2 U1029 ( .A(x_z2[10]), .Z(n1688) );
  HS65_GS_IVX2 U1030 ( .A(x_z2[9]), .Z(n1687) );
  HS65_GS_IVX2 U1031 ( .A(x_z2[8]), .Z(n1686) );
  HS65_GS_IVX2 U1032 ( .A(x_z2[7]), .Z(n1685) );
  HS65_GS_IVX2 U1033 ( .A(x_z2[6]), .Z(n1684) );
  HS65_GS_IVX2 U1034 ( .A(x_z2[5]), .Z(n1683) );
  HS65_GS_IVX2 U1035 ( .A(x_z2[4]), .Z(n1682) );
  HS65_GS_IVX2 U1036 ( .A(x_z2[3]), .Z(n1681) );
  HS65_GS_IVX2 U1037 ( .A(x_z2[2]), .Z(n1680) );
  HS65_GS_IVX2 U1038 ( .A(\mul_b1/fa1_s0[1] ), .Z(n1679) );
  HS65_GS_IVX2 U1039 ( .A(\mul_b1/fa1_s0[0] ), .Z(n1678) );
  HS65_GS_IVX2 U1040 ( .A(n930), .Z(n1378) );
  HS65_GS_HA1X4 U1041 ( .A0(n1679), .B0(n1678), .CO(n1350), .S0(n1652) );
  HS65_GSS_XOR2X3 U1042 ( .A(x_z2[3]), .B(n1652), .Z(\mul_b1/fa1_s0[3] ) );
  HS65_GS_FA1X4 U1043 ( .A0(n933), .B0(n932), .CI(n931), .CO(n940), .S0(n947)
         );
  HS65_GS_FA1X4 U1044 ( .A0(n936), .B0(n935), .CI(n934), .CO(n931), .S0(n946)
         );
  HS65_GS_FA1X4 U1045 ( .A0(n939), .B0(n938), .CI(n937), .CO(n934), .S0(n945)
         );
  HS65_GS_NOR3X1 U1046 ( .A(n947), .B(n946), .C(n945), .Z(n944) );
  HS65_GS_FA1X4 U1047 ( .A0(n942), .B0(n941), .CI(n940), .CO(n523), .S0(n943)
         );
  HS65_GS_IVX2 U1048 ( .A(n943), .Z(n949) );
  HS65_GS_AOI12X2 U1049 ( .A(n944), .B(n949), .C(\mul_b2/result_sat[15] ), .Z(
        n1404) );
  HS65_GS_IVX2 U1050 ( .A(n1404), .Z(n1001) );
  HS65_GS_NAND3X2 U1051 ( .A(n947), .B(n946), .C(n945), .Z(n948) );
  HS65_GS_OAI21X2 U1052 ( .A(n949), .B(n948), .C(\mul_b2/result_sat[15] ), .Z(
        n1405) );
  HS65_GS_IVX2 U1053 ( .A(n1405), .Z(n1397) );
  HS65_GS_AO112X4 U1054 ( .A(n952), .B(n951), .C(n1397), .D(n950), .Z(n953) );
  HS65_GS_NAND2X2 U1055 ( .A(n1001), .B(n953), .Z(\mul_b2/result_sat[0] ) );
  HS65_GS_AO112X4 U1056 ( .A(n956), .B(n955), .C(n1397), .D(n954), .Z(n957) );
  HS65_GS_NAND2X2 U1057 ( .A(n1001), .B(n957), .Z(\mul_b2/result_sat[1] ) );
  HS65_GS_AOI12X2 U1058 ( .A(n960), .B(n959), .C(n1404), .Z(n958) );
  HS65_GS_CBI4I6X2 U1059 ( .A(n960), .B(n959), .C(n958), .D(n1397), .Z(
        \mul_b2/result_sat[2] ) );
  HS65_GS_AO112X4 U1060 ( .A(n963), .B(n962), .C(n1397), .D(n961), .Z(n964) );
  HS65_GS_NAND2X2 U1061 ( .A(n1001), .B(n964), .Z(\mul_b2/result_sat[3] ) );
  HS65_GS_AO112X4 U1062 ( .A(n967), .B(n966), .C(n1397), .D(n965), .Z(n968) );
  HS65_GS_NAND2X2 U1063 ( .A(n1001), .B(n968), .Z(\mul_b2/result_sat[4] ) );
  HS65_GS_AO112X4 U1064 ( .A(n971), .B(n970), .C(n1397), .D(n969), .Z(n972) );
  HS65_GS_NAND2X2 U1065 ( .A(n1001), .B(n972), .Z(\mul_b2/result_sat[5] ) );
  HS65_GS_AO112X4 U1066 ( .A(n975), .B(n974), .C(n1397), .D(n973), .Z(n976) );
  HS65_GS_NAND2X2 U1067 ( .A(n1001), .B(n976), .Z(\mul_b2/result_sat[6] ) );
  HS65_GS_AO112X4 U1068 ( .A(n979), .B(n978), .C(n1397), .D(n977), .Z(n980) );
  HS65_GS_NAND2X2 U1069 ( .A(n1001), .B(n980), .Z(\mul_b2/result_sat[7] ) );
  HS65_GS_AO112X4 U1070 ( .A(n983), .B(n982), .C(n1397), .D(n981), .Z(n984) );
  HS65_GS_NAND2X2 U1071 ( .A(n1001), .B(n984), .Z(\mul_b2/result_sat[8] ) );
  HS65_GS_AO112X4 U1072 ( .A(n987), .B(n986), .C(n1397), .D(n985), .Z(n988) );
  HS65_GS_NAND2X2 U1073 ( .A(n1001), .B(n988), .Z(\mul_b2/result_sat[9] ) );
  HS65_GS_AO112X4 U1074 ( .A(n991), .B(n990), .C(n1397), .D(n989), .Z(n992) );
  HS65_GS_NAND2X2 U1075 ( .A(n1001), .B(n992), .Z(\mul_b2/result_sat[10] ) );
  HS65_GS_AO112X4 U1076 ( .A(n995), .B(n994), .C(n1397), .D(n993), .Z(n996) );
  HS65_GS_NAND2X2 U1077 ( .A(n1001), .B(n996), .Z(\mul_b2/result_sat[11] ) );
  HS65_GS_AO112X4 U1078 ( .A(n999), .B(n998), .C(n1397), .D(n997), .Z(n1000)
         );
  HS65_GS_NAND2X2 U1079 ( .A(n1001), .B(n1000), .Z(\mul_b2/result_sat[12] ) );
  HS65_GS_IVX2 U1080 ( .A(x_reg2[15]), .Z(n1002) );
  HS65_GS_IVX4 U1081 ( .A(n1002), .Z(n1711) );
  HS65_GSS_XNOR2X3 U1082 ( .A(n1004), .B(n1003), .Z(n1020) );
  HS65_GS_NAND2X2 U1083 ( .A(n1007), .B(n1006), .Z(n1005) );
  HS65_GS_OAI21X2 U1084 ( .A(n1007), .B(n1006), .C(n1005), .Z(n1008) );
  HS65_GSS_XOR2X3 U1085 ( .A(n1009), .B(n1008), .Z(n1019) );
  HS65_GS_FA1X4 U1086 ( .A0(n1012), .B0(n1011), .CI(n1010), .CO(n1009), .S0(
        n1018) );
  HS65_GS_FA1X4 U1087 ( .A0(n1015), .B0(n1014), .CI(n1013), .CO(n1010), .S0(
        n1017) );
  HS65_GS_NOR3AX2 U1088 ( .A(n1019), .B(n1018), .C(n1017), .Z(n1016) );
  HS65_GS_AOI12X2 U1089 ( .A(n1020), .B(n1016), .C(\mul_a1/result_sat[15] ), 
        .Z(n1443) );
  HS65_GS_IVX2 U1090 ( .A(n1443), .Z(n1045) );
  HS65_GS_NAND4ABX3 U1091 ( .A(n1020), .B(n1019), .C(n1018), .D(n1017), .Z(
        n1021) );
  HS65_GS_NAND2X2 U1092 ( .A(\mul_a1/result_sat[15] ), .B(n1021), .Z(n1444) );
  HS65_GS_IVX2 U1093 ( .A(n1444), .Z(n1436) );
  HS65_GS_AO112X4 U1094 ( .A(n1024), .B(n1023), .C(n1436), .D(n1022), .Z(n1025) );
  HS65_GS_NAND2X2 U1095 ( .A(n1045), .B(n1025), .Z(\mul_a1/result_sat[0] ) );
  HS65_GSS_XOR2X3 U1096 ( .A(n1027), .B(n1026), .Z(n1030) );
  HS65_GS_OAI21X2 U1097 ( .A(n1029), .B(n1030), .C(n1444), .Z(n1028) );
  HS65_GS_CBI4I1X3 U1098 ( .A(n1030), .B(n1029), .C(n1028), .D(n1045), .Z(
        \mul_a1/result_sat[8] ) );
  HS65_GS_OAI21X2 U1099 ( .A(n1032), .B(n1033), .C(n1444), .Z(n1031) );
  HS65_GS_CBI4I1X3 U1100 ( .A(n1033), .B(n1032), .C(n1031), .D(n1045), .Z(
        \mul_a1/result_sat[9] ) );
  HS65_GS_OAI21X2 U1101 ( .A(n1035), .B(n1036), .C(n1444), .Z(n1034) );
  HS65_GS_CBI4I1X3 U1102 ( .A(n1036), .B(n1035), .C(n1034), .D(n1045), .Z(
        \mul_a1/result_sat[10] ) );
  HS65_GS_AO112X4 U1103 ( .A(n1039), .B(n1038), .C(n1436), .D(n1037), .Z(n1040) );
  HS65_GS_NAND2X2 U1104 ( .A(n1045), .B(n1040), .Z(\mul_a1/result_sat[11] ) );
  HS65_GS_AO112X4 U1105 ( .A(n1043), .B(n1042), .C(n1436), .D(n1041), .Z(n1044) );
  HS65_GS_NAND2X2 U1106 ( .A(n1045), .B(n1044), .Z(\mul_a1/result_sat[12] ) );
  HS65_GS_HA1X4 U1107 ( .A0(n1663), .B0(n1046), .CO(n1472), .S0(n1494) );
  HS65_GS_IVX2 U1108 ( .A(n1494), .Z(n1048) );
  HS65_GS_NAND2X2 U1109 ( .A(n1494), .B(y_z1[12]), .Z(n1047) );
  HS65_GS_CBI4I1X3 U1110 ( .A(n1659), .B(n1048), .C(n1667), .D(n1047), .Z(
        \mul_a1/fa1_c1[18] ) );
  HS65_GS_HA1X4 U1111 ( .A0(n1659), .B0(n1049), .CO(n1475), .S0(n1496) );
  HS65_GS_IVX2 U1112 ( .A(n1496), .Z(n1051) );
  HS65_GS_NAND2X2 U1113 ( .A(n1496), .B(y_z1[14]), .Z(n1050) );
  HS65_GS_CBI4I1X3 U1114 ( .A(n1655), .B(n1051), .C(n1663), .D(n1050), .Z(
        \mul_a1/fa1_c1[20] ) );
  HS65_GS_HA1X4 U1115 ( .A0(n1447), .B0(n1446), .CO(n1052) );
  HS65_GS_HA1X4 U1116 ( .A0(n1484), .B0(n1052), .CO(n1676) );
  HS65_GS_IVX2 U1117 ( .A(n1053), .Z(n1055) );
  HS65_GS_AOI22X1 U1118 ( .A(n1056), .B(n1055), .C(n1057), .D(n1054), .Z(n1071) );
  HS65_GS_AOI12X2 U1119 ( .A(n1059), .B(n1058), .C(n1057), .Z(n1069) );
  HS65_GS_FA1X4 U1120 ( .A0(n1062), .B0(n1061), .CI(n1060), .CO(n732), .S0(
        n1068) );
  HS65_GS_FA1X4 U1121 ( .A0(n1065), .B0(n1064), .CI(n1063), .CO(n1060), .S0(
        n1067) );
  HS65_GS_NOR3X1 U1122 ( .A(n1069), .B(n1068), .C(n1067), .Z(n1066) );
  HS65_GS_AOI12X2 U1123 ( .A(n1071), .B(n1066), .C(\mul_b0/result_sat[15] ), 
        .Z(n1509) );
  HS65_GS_IVX2 U1124 ( .A(n1509), .Z(n1122) );
  HS65_GS_NAND3X2 U1125 ( .A(n1069), .B(n1068), .C(n1067), .Z(n1070) );
  HS65_GS_OAI21X2 U1126 ( .A(n1071), .B(n1070), .C(\mul_b0/result_sat[15] ), 
        .Z(n1510) );
  HS65_GS_IVX2 U1127 ( .A(n1510), .Z(n1502) );
  HS65_GS_AO112X4 U1128 ( .A(n1074), .B(n1073), .C(n1502), .D(n1072), .Z(n1075) );
  HS65_GS_NAND2X2 U1129 ( .A(n1122), .B(n1075), .Z(\mul_b0/result_sat[0] ) );
  HS65_GS_AOI12X2 U1130 ( .A(n1078), .B(n1077), .C(n1509), .Z(n1076) );
  HS65_GS_CBI4I6X2 U1131 ( .A(n1078), .B(n1077), .C(n1076), .D(n1502), .Z(
        \mul_b0/result_sat[1] ) );
  HS65_GS_AO112X4 U1132 ( .A(n1081), .B(n1080), .C(n1502), .D(n1079), .Z(n1082) );
  HS65_GS_NAND2X2 U1133 ( .A(n1122), .B(n1082), .Z(\mul_b0/result_sat[2] ) );
  HS65_GS_AO112X4 U1134 ( .A(n1085), .B(n1084), .C(n1502), .D(n1083), .Z(n1086) );
  HS65_GS_NAND2X2 U1135 ( .A(n1122), .B(n1086), .Z(\mul_b0/result_sat[3] ) );
  HS65_GS_AOI12X2 U1136 ( .A(n1089), .B(n1088), .C(n1509), .Z(n1087) );
  HS65_GS_CBI4I6X2 U1137 ( .A(n1089), .B(n1088), .C(n1087), .D(n1502), .Z(
        \mul_b0/result_sat[4] ) );
  HS65_GS_AO112X4 U1138 ( .A(n1092), .B(n1091), .C(n1502), .D(n1090), .Z(n1093) );
  HS65_GS_NAND2X2 U1139 ( .A(n1122), .B(n1093), .Z(\mul_b0/result_sat[5] ) );
  HS65_GS_AO112X4 U1140 ( .A(n1096), .B(n1095), .C(n1502), .D(n1094), .Z(n1097) );
  HS65_GS_NAND2X2 U1141 ( .A(n1122), .B(n1097), .Z(\mul_b0/result_sat[6] ) );
  HS65_GS_AO112X4 U1142 ( .A(n1100), .B(n1099), .C(n1502), .D(n1098), .Z(n1101) );
  HS65_GS_NAND2X2 U1143 ( .A(n1122), .B(n1101), .Z(\mul_b0/result_sat[7] ) );
  HS65_GS_AO112X4 U1144 ( .A(n1104), .B(n1103), .C(n1502), .D(n1102), .Z(n1105) );
  HS65_GS_NAND2X2 U1145 ( .A(n1122), .B(n1105), .Z(\mul_b0/result_sat[8] ) );
  HS65_GS_AO112X4 U1146 ( .A(n1108), .B(n1107), .C(n1502), .D(n1106), .Z(n1109) );
  HS65_GS_NAND2X2 U1147 ( .A(n1122), .B(n1109), .Z(\mul_b0/result_sat[9] ) );
  HS65_GS_AO112X4 U1148 ( .A(n1112), .B(n1111), .C(n1502), .D(n1110), .Z(n1113) );
  HS65_GS_NAND2X2 U1149 ( .A(n1122), .B(n1113), .Z(\mul_b0/result_sat[10] ) );
  HS65_GS_AO112X4 U1150 ( .A(n1116), .B(n1115), .C(n1502), .D(n1114), .Z(n1117) );
  HS65_GS_NAND2X2 U1151 ( .A(n1122), .B(n1117), .Z(\mul_b0/result_sat[11] ) );
  HS65_GS_AO112X4 U1152 ( .A(n1120), .B(n1119), .C(n1502), .D(n1118), .Z(n1121) );
  HS65_GS_NAND2X2 U1153 ( .A(n1122), .B(n1121), .Z(\mul_b0/result_sat[12] ) );
  HS65_GS_IVX2 U1154 ( .A(n1554), .Z(n1713) );
  HS65_GSS_XOR2X3 U1155 ( .A(n1124), .B(n1123), .Z(n1145) );
  HS65_GS_FA1X4 U1156 ( .A0(n1127), .B0(n1126), .CI(n1125), .CO(n1130), .S0(
        n1128) );
  HS65_GS_IVX2 U1157 ( .A(n1128), .Z(n1143) );
  HS65_GS_FA1X4 U1158 ( .A0(n1131), .B0(n1130), .CI(n1129), .CO(n1136), .S0(
        n1141) );
  HS65_GS_FA1X4 U1159 ( .A0(n1134), .B0(n1133), .CI(n1132), .CO(n1126), .S0(
        n1140) );
  HS65_GS_FA1X4 U1160 ( .A0(n1137), .B0(n1136), .CI(n1135), .CO(n198), .S0(
        n1139) );
  HS65_GS_NAND3X2 U1161 ( .A(n1141), .B(n1140), .C(n1139), .Z(n1138) );
  HS65_GS_OAI12X3 U1162 ( .A(n1143), .B(n1138), .C(\mul_b1/result_sat[15] ), 
        .Z(n1607) );
  HS65_GS_OAI21X2 U1163 ( .A(n1145), .B(n1146), .C(n1607), .Z(n1144) );
  HS65_GS_NOR3X1 U1164 ( .A(n1141), .B(n1140), .C(n1139), .Z(n1142) );
  HS65_GS_AOI12X3 U1165 ( .A(n1143), .B(n1142), .C(\mul_b1/result_sat[15] ), 
        .Z(n1609) );
  HS65_GS_IVX2 U1166 ( .A(n1609), .Z(n1150) );
  HS65_GS_CBI4I1X3 U1167 ( .A(n1146), .B(n1145), .C(n1144), .D(n1150), .Z(
        \mul_b1/result_sat[0] ) );
  HS65_GS_AOI12X2 U1168 ( .A(n1149), .B(n1148), .C(n1147), .Z(n1152) );
  HS65_GS_OAI21X2 U1169 ( .A(n1152), .B(n1153), .C(n1607), .Z(n1151) );
  HS65_GS_CBI4I1X3 U1170 ( .A(n1153), .B(n1152), .C(n1151), .D(n1150), .Z(
        \mul_b1/result_sat[7] ) );
  HS65_GS_IVX2 U1171 ( .A(n1693), .Z(n1712) );
  HS65_GS_NOR2X2 U1172 ( .A(n1678), .B(n1680), .Z(\mul_b1/fa1_c1[8] ) );
  HS65_GS_NOR2X2 U1173 ( .A(n1679), .B(n1681), .Z(\mul_b1/fa1_c1[9] ) );
  HS65_GS_NOR2X2 U1174 ( .A(n1680), .B(n1682), .Z(\mul_b1/fa1_c1[10] ) );
  HS65_GS_NOR2X2 U1175 ( .A(n1681), .B(n1683), .Z(\mul_b1/fa1_c1[11] ) );
  HS65_GS_NOR2X2 U1176 ( .A(n1682), .B(n1684), .Z(\mul_b1/fa1_c1[12] ) );
  HS65_GS_NOR2X2 U1177 ( .A(n1683), .B(n1685), .Z(\mul_b1/fa1_c1[13] ) );
  HS65_GS_NOR2X2 U1178 ( .A(n1684), .B(n1686), .Z(\mul_b1/fa1_c1[14] ) );
  HS65_GS_NOR2X2 U1179 ( .A(n1685), .B(n1687), .Z(\mul_b1/fa1_c1[15] ) );
  HS65_GS_NOR2X2 U1180 ( .A(n1686), .B(n1688), .Z(\mul_b1/fa1_c1[16] ) );
  HS65_GS_NOR2X2 U1181 ( .A(n1687), .B(n1689), .Z(\mul_b1/fa1_c1[17] ) );
  HS65_GS_NOR2X2 U1182 ( .A(n1688), .B(n1690), .Z(\mul_b1/fa1_c1[18] ) );
  HS65_GS_NOR2X2 U1183 ( .A(n1689), .B(n1691), .Z(\mul_b1/fa1_c1[19] ) );
  HS65_GS_NOR2X2 U1184 ( .A(n1690), .B(n1692), .Z(\mul_b1/fa1_c1[20] ) );
  HS65_GS_NOR2X2 U1185 ( .A(n1693), .B(n1691), .Z(\mul_b1/fa1_c1[21] ) );
  HS65_GS_NOR2X2 U1186 ( .A(n1693), .B(n1692), .Z(\mul_b1/fa1_c1[22] ) );
  HS65_GS_IVX2 U1187 ( .A(x_z1[14]), .Z(n1548) );
  HS65_GS_IVX2 U1188 ( .A(x_z1[13]), .Z(n1546) );
  HS65_GS_IVX2 U1189 ( .A(x_z1[12]), .Z(n1544) );
  HS65_GS_IVX2 U1190 ( .A(x_z1[11]), .Z(n1542) );
  HS65_GS_IVX2 U1191 ( .A(x_z1[10]), .Z(n1540) );
  HS65_GS_IVX2 U1192 ( .A(x_z1[9]), .Z(n1538) );
  HS65_GS_IVX2 U1193 ( .A(x_z1[8]), .Z(n1536) );
  HS65_GS_IVX2 U1194 ( .A(x_z1[7]), .Z(n1534) );
  HS65_GS_IVX2 U1195 ( .A(x_z1[6]), .Z(n1532) );
  HS65_GS_IVX2 U1196 ( .A(x_z1[5]), .Z(n1521) );
  HS65_GS_IVX2 U1197 ( .A(x_z1[4]), .Z(n1519) );
  HS65_GS_IVX2 U1198 ( .A(x_z1[3]), .Z(n1517) );
  HS65_GS_IVX2 U1199 ( .A(x_z1[2]), .Z(n1515) );
  HS65_GS_IVX2 U1200 ( .A(x_z1[1]), .Z(n1513) );
  HS65_GS_IVX2 U1201 ( .A(x_z1[0]), .Z(n1512) );
  HS65_GSS_XNOR2X3 U1202 ( .A(x_z1[15]), .B(n1154), .Z(n1531) );
  HS65_GSS_XNOR2X3 U1203 ( .A(n1531), .B(n1554), .Z(\mul_b0/fa1_s0[20] ) );
  HS65_GS_NOR2X2 U1204 ( .A(x_z1[15]), .B(n1154), .Z(n1155) );
  HS65_GSS_XNOR2X3 U1205 ( .A(n1155), .B(n1554), .Z(\mul_b0/fa1_s0[31] ) );
  HS65_GS_HA1X4 U1206 ( .A0(n1317), .B0(n1247), .CO(n1170), .S0(n1218) );
  HS65_GSS_XOR2X3 U1207 ( .A(n1218), .B(y_z2[0]), .Z(\mul_a2/fa1_s1[10] ) );
  HS65_GS_HA1X4 U1208 ( .A0(n1331), .B0(n1156), .CO(n1172), .S0(n1234) );
  HS65_GS_HA1X4 U1209 ( .A0(n1333), .B0(n1157), .CO(n1171), .S0(n1233) );
  HS65_GSS_XOR2X3 U1210 ( .A(n1234), .B(n1233), .Z(\mul_a2/fa1_s1[18] ) );
  HS65_GS_HA1X4 U1211 ( .A0(n1329), .B0(n1158), .CO(n1156), .S0(n1232) );
  HS65_GS_HA1X4 U1212 ( .A0(n1331), .B0(n1159), .CO(n1157), .S0(n1231) );
  HS65_GSS_XOR2X3 U1213 ( .A(n1232), .B(n1231), .Z(\mul_a2/fa1_s1[17] ) );
  HS65_GS_HA1X4 U1214 ( .A0(n1329), .B0(n1160), .CO(n1159), .S0(n1230) );
  HS65_GS_HA1X4 U1215 ( .A0(n1327), .B0(n1161), .CO(n1158), .S0(n1229) );
  HS65_GSS_XOR2X3 U1216 ( .A(n1230), .B(n1229), .Z(\mul_a2/fa1_s1[16] ) );
  HS65_GS_HA1X4 U1217 ( .A0(n1325), .B0(n1162), .CO(n1161), .S0(n1228) );
  HS65_GS_HA1X4 U1218 ( .A0(n1327), .B0(n1163), .CO(n1160), .S0(n1227) );
  HS65_GSS_XOR2X3 U1219 ( .A(n1228), .B(n1227), .Z(\mul_a2/fa1_s1[15] ) );
  HS65_GS_HA1X4 U1220 ( .A0(n1323), .B0(n1164), .CO(n1162), .S0(n1226) );
  HS65_GS_HA1X4 U1221 ( .A0(n1325), .B0(n1165), .CO(n1163), .S0(n1225) );
  HS65_GSS_XOR2X3 U1222 ( .A(n1226), .B(n1225), .Z(\mul_a2/fa1_s1[14] ) );
  HS65_GS_HA1X4 U1223 ( .A0(n1321), .B0(n1166), .CO(n1164), .S0(n1224) );
  HS65_GS_HA1X4 U1224 ( .A0(n1323), .B0(n1167), .CO(n1165), .S0(n1223) );
  HS65_GSS_XOR2X3 U1225 ( .A(n1224), .B(n1223), .Z(\mul_a2/fa1_s1[13] ) );
  HS65_GS_HA1X4 U1226 ( .A0(n1321), .B0(n1168), .CO(n1167), .S0(n1222) );
  HS65_GS_HA1X4 U1227 ( .A0(n1319), .B0(n1169), .CO(n1166), .S0(n1221) );
  HS65_GSS_XOR2X3 U1228 ( .A(n1222), .B(n1221), .Z(\mul_a2/fa1_s1[12] ) );
  HS65_GS_HA1X4 U1229 ( .A0(n1319), .B0(n1170), .CO(n1168), .S0(n1220) );
  HS65_GS_HA1X4 U1230 ( .A0(n1317), .B0(n1247), .CO(n1169), .S0(n1219) );
  HS65_GSS_XOR2X3 U1231 ( .A(n1220), .B(n1219), .Z(\mul_a2/fa1_s1[11] ) );
  HS65_GS_AND2X4 U1232 ( .A(n1322), .B(y_z2[3]), .Z(\mul_a2/fa1_c0[5] ) );
  HS65_GS_HA1X4 U1233 ( .A0(n1335), .B0(n1171), .CO(n1174), .S0(n1236) );
  HS65_GS_HA1X4 U1234 ( .A0(n1333), .B0(n1172), .CO(n1173), .S0(n1235) );
  HS65_GSS_XOR2X3 U1235 ( .A(n1236), .B(n1235), .Z(\mul_a2/fa1_s1[19] ) );
  HS65_GS_HA1X4 U1236 ( .A0(n1335), .B0(n1173), .CO(n1175), .S0(n1238) );
  HS65_GS_HA1X4 U1237 ( .A0(n1337), .B0(n1174), .CO(n1176), .S0(n1237) );
  HS65_GSS_XOR2X3 U1238 ( .A(n1238), .B(n1237), .Z(\mul_a2/fa1_s1[20] ) );
  HS65_GS_HA1X4 U1239 ( .A0(n1337), .B0(n1175), .CO(n1177), .S0(n1240) );
  HS65_GS_HA1X4 U1240 ( .A0(n1339), .B0(n1176), .CO(n1178), .S0(n1239) );
  HS65_GSS_XOR2X3 U1241 ( .A(n1240), .B(n1239), .Z(\mul_a2/fa1_s1[21] ) );
  HS65_GS_HA1X4 U1242 ( .A0(n1339), .B0(n1177), .CO(n1180), .S0(n1242) );
  HS65_GS_HA1X4 U1243 ( .A0(n1341), .B0(n1178), .CO(n1179), .S0(n1241) );
  HS65_GSS_XOR2X3 U1244 ( .A(n1242), .B(n1241), .Z(\mul_a2/fa1_s1[22] ) );
  HS65_GS_HA1X4 U1245 ( .A0(n1343), .B0(n1179), .CO(n1182), .S0(n1244) );
  HS65_GS_HA1X4 U1246 ( .A0(n1341), .B0(n1180), .CO(n1181), .S0(n1243) );
  HS65_GSS_XOR2X3 U1247 ( .A(n1244), .B(n1243), .Z(\mul_a2/fa1_s1[23] ) );
  HS65_GS_HA1X4 U1248 ( .A0(n1343), .B0(n1181), .CO(n871), .S0(n1246) );
  HS65_GSS_XNOR2X3 U1249 ( .A(y_z2[15]), .B(n1182), .Z(n1245) );
  HS65_GSS_XOR2X3 U1250 ( .A(n1246), .B(n1245), .Z(\mul_a2/fa1_s1[24] ) );
  HS65_GS_HA1X4 U1251 ( .A0(n1317), .B0(n1247), .CO(n1184), .S0(n1183) );
  HS65_GS_AND2X4 U1252 ( .A(y_z2[0]), .B(n1183), .Z(\mul_a2/fa1_c0[2] ) );
  HS65_GS_HA1X4 U1253 ( .A0(n1319), .B0(n1184), .CO(n1185), .S0(n1318) );
  HS65_GS_AND2X4 U1254 ( .A(n1318), .B(y_z2[1]), .Z(\mul_a2/fa1_c0[3] ) );
  HS65_GS_HA1X4 U1255 ( .A0(n1321), .B0(n1185), .CO(n1186), .S0(n1320) );
  HS65_GS_AND2X4 U1256 ( .A(n1320), .B(y_z2[2]), .Z(\mul_a2/fa1_c0[4] ) );
  HS65_GS_HA1X4 U1257 ( .A0(n1323), .B0(n1186), .CO(n1307), .S0(n1322) );
  HS65_GS_AND2X4 U1258 ( .A(n1324), .B(y_z2[4]), .Z(\mul_a2/fa1_c0[6] ) );
  HS65_GS_IVX2 U1259 ( .A(n1216), .Z(n1701) );
  HS65_GS_OAI21X2 U1260 ( .A(n1189), .B(n1188), .C(n1187), .Z(n1190) );
  HS65_GS_OAI21X2 U1261 ( .A(n1701), .B(n1190), .C(n1702), .Z(
        \mul_a2/result_sat[0] ) );
  HS65_GS_OAI21X2 U1262 ( .A(n1193), .B(n1192), .C(n1191), .Z(n1194) );
  HS65_GS_OAI21X2 U1263 ( .A(n1701), .B(n1194), .C(n1702), .Z(
        \mul_a2/result_sat[1] ) );
  HS65_GS_OAI21X2 U1264 ( .A(n1197), .B(n1196), .C(n1195), .Z(n1198) );
  HS65_GS_OAI21X2 U1265 ( .A(n1701), .B(n1198), .C(n1702), .Z(
        \mul_a2/result_sat[3] ) );
  HS65_GSS_XOR2X3 U1266 ( .A(n1200), .B(n1199), .Z(n1201) );
  HS65_GSS_XNOR2X3 U1267 ( .A(n1202), .B(n1201), .Z(n1203) );
  HS65_GS_OAI21X2 U1268 ( .A(n1701), .B(n1203), .C(n1702), .Z(
        \mul_a2/result_sat[4] ) );
  HS65_GS_OAI21X2 U1269 ( .A(n1206), .B(n1205), .C(n1204), .Z(n1207) );
  HS65_GS_OAI21X2 U1270 ( .A(n1701), .B(n1207), .C(n1702), .Z(
        \mul_a2/result_sat[6] ) );
  HS65_GS_FA1X4 U1271 ( .A0(n1210), .B0(n1209), .CI(n1208), .CO(n1212), .S0(
        n1211) );
  HS65_GS_OA12X4 U1272 ( .A(n1215), .B(n1211), .C(n1216), .Z(
        \mul_a2/result_sat[10] ) );
  HS65_GS_FA1X4 U1273 ( .A0(n1214), .B0(n1213), .CI(n1212), .CO(n917), .S0(
        n1217) );
  HS65_GS_AO12X4 U1274 ( .A(n1217), .B(n1216), .C(n1215), .Z(
        \mul_a2/result_sat[11] ) );
  HS65_GS_AND2X4 U1275 ( .A(n1218), .B(y_z2[0]), .Z(\mul_a2/fa1_c1[10] ) );
  HS65_GS_AND2X4 U1276 ( .A(n1220), .B(n1219), .Z(\mul_a2/fa1_c1[11] ) );
  HS65_GS_AND2X4 U1277 ( .A(n1222), .B(n1221), .Z(\mul_a2/fa1_c1[12] ) );
  HS65_GS_AND2X4 U1278 ( .A(n1224), .B(n1223), .Z(\mul_a2/fa1_c1[13] ) );
  HS65_GS_AND2X4 U1279 ( .A(n1226), .B(n1225), .Z(\mul_a2/fa1_c1[14] ) );
  HS65_GS_AND2X4 U1280 ( .A(n1228), .B(n1227), .Z(\mul_a2/fa1_c1[15] ) );
  HS65_GS_AND2X4 U1281 ( .A(n1230), .B(n1229), .Z(\mul_a2/fa1_c1[16] ) );
  HS65_GS_AND2X4 U1282 ( .A(n1232), .B(n1231), .Z(\mul_a2/fa1_c1[17] ) );
  HS65_GS_AND2X4 U1283 ( .A(n1234), .B(n1233), .Z(\mul_a2/fa1_c1[18] ) );
  HS65_GS_AND2X4 U1284 ( .A(n1236), .B(n1235), .Z(\mul_a2/fa1_c1[19] ) );
  HS65_GS_AND2X4 U1285 ( .A(n1238), .B(n1237), .Z(\mul_a2/fa1_c1[20] ) );
  HS65_GS_AND2X4 U1286 ( .A(n1240), .B(n1239), .Z(\mul_a2/fa1_c1[21] ) );
  HS65_GS_AND2X4 U1287 ( .A(n1242), .B(n1241), .Z(\mul_a2/fa1_c1[22] ) );
  HS65_GS_AND2X4 U1288 ( .A(n1244), .B(n1243), .Z(\mul_a2/fa1_c1[23] ) );
  HS65_GS_AND2X4 U1289 ( .A(n1246), .B(n1245), .Z(\mul_a2/fa1_c1[24] ) );
  HS65_GS_MUX21X4 U1290 ( .D0(n1713), .D1(data_in[15]), .S0(valid_in), .Z(
        n1715) );
  HS65_GS_MUX21X4 U1291 ( .D0(x_z1[14]), .D1(data_in[14]), .S0(valid_in), .Z(
        n1716) );
  HS65_GS_MUX21X4 U1292 ( .D0(x_z1[13]), .D1(data_in[13]), .S0(n1714), .Z(
        n1717) );
  HS65_GS_MUX21X4 U1293 ( .D0(x_z1[12]), .D1(data_in[12]), .S0(valid_in), .Z(
        n1718) );
  HS65_GS_BFX4 U1294 ( .A(valid_in), .Z(n1306) );
  HS65_GS_MUX21X4 U1295 ( .D0(x_z1[11]), .D1(data_in[11]), .S0(n1306), .Z(
        n1719) );
  HS65_GS_MUX21X4 U1296 ( .D0(x_z1[10]), .D1(data_in[10]), .S0(n1714), .Z(
        n1720) );
  HS65_GS_MUX21X4 U1297 ( .D0(x_z1[9]), .D1(data_in[9]), .S0(valid_in), .Z(
        n1721) );
  HS65_GS_MUX21X4 U1298 ( .D0(x_z1[8]), .D1(data_in[8]), .S0(n1305), .Z(n1722)
         );
  HS65_GS_MUX21X4 U1299 ( .D0(x_z1[7]), .D1(data_in[7]), .S0(n1714), .Z(n1723)
         );
  HS65_GS_MUX21X4 U1300 ( .D0(x_z1[6]), .D1(data_in[6]), .S0(n1714), .Z(n1724)
         );
  HS65_GS_MUX21X4 U1301 ( .D0(x_z1[5]), .D1(data_in[5]), .S0(n1714), .Z(n1725)
         );
  HS65_GS_MUX21X4 U1302 ( .D0(x_z1[4]), .D1(data_in[4]), .S0(n1714), .Z(n1726)
         );
  HS65_GS_MUX21X4 U1303 ( .D0(x_z1[3]), .D1(data_in[3]), .S0(n1714), .Z(n1727)
         );
  HS65_GS_MUXI21X2 U1304 ( .D0(n1247), .D1(n1446), .S0(n1306), .Z(n1810) );
  HS65_GS_MUX21X4 U1305 ( .D0(x_z1[2]), .D1(data_in[2]), .S0(n1714), .Z(n1728)
         );
  HS65_GS_MUX21X4 U1306 ( .D0(x_z1[1]), .D1(data_in[1]), .S0(n1714), .Z(n1729)
         );
  HS65_GS_MUXI21X2 U1307 ( .D0(n1317), .D1(n1447), .S0(n1290), .Z(n1807) );
  HS65_GS_MUX21X4 U1308 ( .D0(x_z1[0]), .D1(data_in[0]), .S0(valid_in), .Z(
        n1730) );
  HS65_GS_MUXI21X2 U1309 ( .D0(n1693), .D1(n1554), .S0(n1306), .Z(n1731) );
  HS65_GS_OAI112X1 U1310 ( .A(n1249), .B(p_a1[1]), .C(n1291), .D(n1248), .Z(
        n1250) );
  HS65_GS_AO22X4 U1311 ( .A(data_out[1]), .B(n1706), .C(n1292), .D(n1250), .Z(
        n1805) );
  HS65_GS_MUXI21X2 U1312 ( .D0(n1002), .D1(n1693), .S0(n1306), .Z(n1732) );
  HS65_GS_MUXI21X2 U1313 ( .D0(n1319), .D1(n1484), .S0(n1290), .Z(n1804) );
  HS65_GS_MUXI21X2 U1314 ( .D0(n1692), .D1(n1548), .S0(n1306), .Z(n1733) );
  HS65_GS_MUX21X4 U1315 ( .D0(x_reg2[14]), .D1(x_z2[14]), .S0(n1714), .Z(n1734) );
  HS65_GS_OAI112X1 U1316 ( .A(n1253), .B(n1252), .C(n1291), .D(n1251), .Z(
        n1254) );
  HS65_GS_AO22X4 U1317 ( .A(data_out[2]), .B(n1706), .C(n1292), .D(n1254), .Z(
        n1802) );
  HS65_GS_MUXI21X2 U1318 ( .D0(n1691), .D1(n1546), .S0(n1306), .Z(n1735) );
  HS65_GS_MUXI21X2 U1319 ( .D0(n1321), .D1(n1677), .S0(n1290), .Z(n1801) );
  HS65_GS_AOI112X2 U1320 ( .A(n1257), .B(n1256), .C(n1304), .D(n1255), .Z(
        n1258) );
  HS65_GS_AO112X4 U1321 ( .A(data_out[3]), .B(n1706), .C(n1258), .D(n1301), 
        .Z(n1799) );
  HS65_GS_MUX21X4 U1322 ( .D0(x_reg2[13]), .D1(x_z2[13]), .S0(n1305), .Z(n1736) );
  HS65_GS_MUXI21X2 U1323 ( .D0(n1323), .D1(n1675), .S0(n1290), .Z(n1798) );
  HS65_GS_OAI112X1 U1324 ( .A(n1261), .B(n1260), .C(n1291), .D(n1259), .Z(
        n1262) );
  HS65_GS_AO22X4 U1325 ( .A(data_out[4]), .B(n1706), .C(n1292), .D(n1262), .Z(
        n1796) );
  HS65_GS_MUXI21X2 U1326 ( .D0(n1690), .D1(n1544), .S0(n1306), .Z(n1737) );
  HS65_GS_MUXI21X2 U1327 ( .D0(n1325), .D1(n1673), .S0(n1306), .Z(n1795) );
  HS65_GS_OAI112X1 U1328 ( .A(n1265), .B(n1264), .C(n1291), .D(n1263), .Z(
        n1266) );
  HS65_GS_AO22X4 U1329 ( .A(data_out[5]), .B(n1706), .C(n1292), .D(n1266), .Z(
        n1793) );
  HS65_GS_MUX21X4 U1330 ( .D0(x_reg2[12]), .D1(x_z2[12]), .S0(valid_in), .Z(
        n1738) );
  HS65_GS_MUXI21X2 U1331 ( .D0(n1327), .D1(n1671), .S0(n1290), .Z(n1792) );
  HS65_GS_OAI112X1 U1332 ( .A(n1269), .B(n1268), .C(n1291), .D(n1267), .Z(
        n1270) );
  HS65_GS_AO22X4 U1333 ( .A(data_out[6]), .B(n1706), .C(n1292), .D(n1270), .Z(
        n1790) );
  HS65_GS_MUXI21X2 U1334 ( .D0(n1329), .D1(n1669), .S0(n1290), .Z(n1789) );
  HS65_GS_MUXI21X2 U1335 ( .D0(n1689), .D1(n1542), .S0(n1305), .Z(n1739) );
  HS65_GS_OAI112X1 U1336 ( .A(n1273), .B(n1272), .C(n1291), .D(n1271), .Z(
        n1274) );
  HS65_GS_AO22X4 U1337 ( .A(data_out[7]), .B(n1706), .C(n1292), .D(n1274), .Z(
        n1787) );
  HS65_GS_MUXI21X2 U1338 ( .D0(n1331), .D1(n1667), .S0(n1290), .Z(n1786) );
  HS65_GS_MUX21X4 U1339 ( .D0(x_reg2[11]), .D1(x_z2[11]), .S0(n1714), .Z(n1740) );
  HS65_GS_OAI112X1 U1340 ( .A(n1277), .B(n1276), .C(n1291), .D(n1275), .Z(
        n1278) );
  HS65_GS_AO22X4 U1341 ( .A(data_out[8]), .B(n1706), .C(n1292), .D(n1278), .Z(
        n1784) );
  HS65_GS_MUXI21X2 U1342 ( .D0(n1688), .D1(n1540), .S0(n1305), .Z(n1741) );
  HS65_GS_MUXI21X2 U1343 ( .D0(n1333), .D1(n1665), .S0(n1290), .Z(n1783) );
  HS65_GS_OAI112X1 U1344 ( .A(n1281), .B(n1280), .C(n1291), .D(n1279), .Z(
        n1282) );
  HS65_GS_AO22X4 U1345 ( .A(data_out[9]), .B(n1706), .C(n1292), .D(n1282), .Z(
        n1781) );
  HS65_GS_MUX21X4 U1346 ( .D0(x_reg2[10]), .D1(x_z2[10]), .S0(n1714), .Z(n1742) );
  HS65_GS_MUXI21X2 U1347 ( .D0(n1335), .D1(n1663), .S0(n1306), .Z(n1780) );
  HS65_GS_MUXI21X2 U1348 ( .D0(n1687), .D1(n1538), .S0(n1305), .Z(n1743) );
  HS65_GS_IVX2 U1349 ( .A(data_out[10]), .Z(n1289) );
  HS65_GS_MUXI21X2 U1350 ( .D0(n1663), .D1(n1289), .S0(n1290), .Z(n1779) );
  HS65_GS_MUX21X4 U1351 ( .D0(x_reg2[9]), .D1(x_z2[9]), .S0(n1306), .Z(n1744)
         );
  HS65_GSS_XOR2X3 U1352 ( .A(n1284), .B(n1283), .Z(n1287) );
  HS65_GS_OAI21X2 U1353 ( .A(n1286), .B(n1287), .C(n1291), .Z(n1285) );
  HS65_GS_CBI4I1X3 U1354 ( .A(n1287), .B(n1286), .C(n1285), .D(n1292), .Z(
        n1288) );
  HS65_GS_OAI21X2 U1355 ( .A(valid_T3), .B(n1289), .C(n1288), .Z(n1778) );
  HS65_GS_MUXI21X2 U1356 ( .D0(n1686), .D1(n1536), .S0(n1305), .Z(n1745) );
  HS65_GS_MUXI21X2 U1357 ( .D0(n1337), .D1(n1661), .S0(n1290), .Z(n1777) );
  HS65_GS_MUX21X4 U1358 ( .D0(x_reg2[8]), .D1(x_z2[8]), .S0(valid_in), .Z(
        n1746) );
  HS65_GS_IVX2 U1359 ( .A(data_out[11]), .Z(n1297) );
  HS65_GS_MUXI21X2 U1360 ( .D0(n1661), .D1(n1297), .S0(n1306), .Z(n1776) );
  HS65_GS_MUXI21X2 U1361 ( .D0(n1685), .D1(n1534), .S0(n1305), .Z(n1747) );
  HS65_GS_OAI21X2 U1362 ( .A(n1294), .B(n1295), .C(n1291), .Z(n1293) );
  HS65_GS_CBI4I1X3 U1363 ( .A(n1295), .B(n1294), .C(n1293), .D(n1292), .Z(
        n1296) );
  HS65_GS_OAI21X2 U1364 ( .A(valid_T3), .B(n1297), .C(n1296), .Z(n1775) );
  HS65_GS_MUX21X4 U1365 ( .D0(x_reg2[7]), .D1(x_z2[7]), .S0(valid_in), .Z(
        n1748) );
  HS65_GS_MUXI21X2 U1366 ( .D0(n1684), .D1(n1532), .S0(n1305), .Z(n1749) );
  HS65_GS_MUX21X4 U1367 ( .D0(x_reg2[6]), .D1(x_z2[6]), .S0(n1306), .Z(n1750)
         );
  HS65_GS_MUXI21X2 U1368 ( .D0(n1683), .D1(n1521), .S0(n1305), .Z(n1751) );
  HS65_GS_MUXI21X2 U1369 ( .D0(n1339), .D1(n1659), .S0(n1306), .Z(n1774) );
  HS65_GS_MUX21X4 U1370 ( .D0(x_reg2[5]), .D1(x_z2[5]), .S0(n1714), .Z(n1752)
         );
  HS65_GS_MUXI21X2 U1371 ( .D0(n1682), .D1(n1519), .S0(n1305), .Z(n1753) );
  HS65_GS_MUX21X4 U1372 ( .D0(x_reg2[4]), .D1(x_z2[4]), .S0(n1306), .Z(n1754)
         );
  HS65_GS_FA1X4 U1373 ( .A0(n1300), .B0(n1299), .CI(n1298), .CO(n926), .S0(
        n1303) );
  HS65_GS_AOI12X2 U1374 ( .A(data_out[12]), .B(n1706), .C(n1301), .Z(n1302) );
  HS65_GS_OAI21X2 U1375 ( .A(n1304), .B(n1303), .C(n1302), .Z(n1772) );
  HS65_GS_MUXI21X2 U1376 ( .D0(n1681), .D1(n1517), .S0(n1305), .Z(n1755) );
  HS65_GS_MUX21X4 U1377 ( .D0(x_reg2[3]), .D1(x_z2[3]), .S0(n1714), .Z(n1756)
         );
  HS65_GS_MUXI21X2 U1378 ( .D0(n1341), .D1(n1657), .S0(n1306), .Z(n1771) );
  HS65_GS_MUXI21X2 U1379 ( .D0(n1680), .D1(n1515), .S0(n1305), .Z(n1757) );
  HS65_GS_MUX21X4 U1380 ( .D0(x_reg2[2]), .D1(x_z2[2]), .S0(valid_in), .Z(
        n1758) );
  HS65_GS_MUXI21X2 U1381 ( .D0(n1679), .D1(n1513), .S0(n1305), .Z(n1759) );
  HS65_GS_MUX21X4 U1382 ( .D0(\mul_b2/fa1_s1[7] ), .D1(\mul_b1/fa1_s0[1] ), 
        .S0(n1714), .Z(n1760) );
  HS65_GS_MUXI21X2 U1383 ( .D0(n1678), .D1(n1512), .S0(n1305), .Z(n1761) );
  HS65_GS_MUX21X4 U1384 ( .D0(x_reg2[0]), .D1(\mul_b1/fa1_s0[0] ), .S0(
        valid_in), .Z(n1762) );
  HS65_GS_IVX2 U1385 ( .A(data_out[15]), .Z(n1705) );
  HS65_GS_MUXI21X2 U1386 ( .D0(n1483), .D1(n1705), .S0(n1306), .Z(n1764) );
  HS65_GS_MUXI21X2 U1387 ( .D0(n1346), .D1(n1483), .S0(n1305), .Z(n1765) );
  HS65_GS_MUXI21X2 U1388 ( .D0(n1343), .D1(n1655), .S0(n1306), .Z(n1768) );
  HS65_GS_HA1X4 U1389 ( .A0(n1325), .B0(n1307), .CO(n1308), .S0(n1324) );
  HS65_GS_AND2X4 U1390 ( .A(n1326), .B(y_z2[5]), .Z(\mul_a2/fa1_c0[7] ) );
  HS65_GS_HA1X4 U1391 ( .A0(n1327), .B0(n1308), .CO(n1309), .S0(n1326) );
  HS65_GS_AND2X4 U1392 ( .A(n1328), .B(y_z2[6]), .Z(\mul_a2/fa1_c0[8] ) );
  HS65_GS_HA1X4 U1393 ( .A0(n1329), .B0(n1309), .CO(n1310), .S0(n1328) );
  HS65_GS_AND2X4 U1394 ( .A(y_z2[7]), .B(n1330), .Z(\mul_a2/fa1_c0[9] ) );
  HS65_GS_HA1X4 U1395 ( .A0(n1331), .B0(n1310), .CO(n1311), .S0(n1330) );
  HS65_GS_AND2X4 U1396 ( .A(n1332), .B(y_z2[8]), .Z(\mul_a2/fa1_c0[10] ) );
  HS65_GS_HA1X4 U1397 ( .A0(n1333), .B0(n1311), .CO(n1312), .S0(n1332) );
  HS65_GS_AND2X4 U1398 ( .A(y_z2[9]), .B(n1334), .Z(\mul_a2/fa1_c0[11] ) );
  HS65_GS_HA1X4 U1399 ( .A0(n1335), .B0(n1312), .CO(n1313), .S0(n1334) );
  HS65_GS_AND2X4 U1400 ( .A(n1336), .B(y_z2[10]), .Z(\mul_a2/fa1_c0[12] ) );
  HS65_GS_HA1X4 U1401 ( .A0(n1337), .B0(n1313), .CO(n1314), .S0(n1336) );
  HS65_GS_AND2X4 U1402 ( .A(n1338), .B(y_z2[11]), .Z(\mul_a2/fa1_c0[13] ) );
  HS65_GS_HA1X4 U1403 ( .A0(n1339), .B0(n1314), .CO(n1315), .S0(n1338) );
  HS65_GS_AND2X4 U1404 ( .A(n1340), .B(y_z2[12]), .Z(\mul_a2/fa1_c0[14] ) );
  HS65_GS_HA1X4 U1405 ( .A0(n1341), .B0(n1315), .CO(n1316), .S0(n1340) );
  HS65_GS_AND2X4 U1406 ( .A(n1342), .B(y_z2[13]), .Z(\mul_a2/fa1_c0[15] ) );
  HS65_GS_HA1X4 U1407 ( .A0(n1343), .B0(n1316), .CO(n1345), .S0(n1342) );
  HS65_GSS_XNOR2X3 U1408 ( .A(y_z2[15]), .B(n1345), .Z(n1344) );
  HS65_GS_AND2X4 U1409 ( .A(y_z2[14]), .B(n1344), .Z(\mul_a2/fa1_c0[16] ) );
  HS65_GSS_XNOR2X3 U1410 ( .A(n1318), .B(n1317), .Z(\mul_a2/fa1_s0[3] ) );
  HS65_GSS_XNOR2X3 U1411 ( .A(n1320), .B(n1319), .Z(\mul_a2/fa1_s0[4] ) );
  HS65_GSS_XNOR2X3 U1412 ( .A(n1322), .B(n1321), .Z(\mul_a2/fa1_s0[5] ) );
  HS65_GSS_XNOR2X3 U1413 ( .A(n1324), .B(n1323), .Z(\mul_a2/fa1_s0[6] ) );
  HS65_GSS_XNOR2X3 U1414 ( .A(n1326), .B(n1325), .Z(\mul_a2/fa1_s0[7] ) );
  HS65_GSS_XNOR2X3 U1415 ( .A(n1328), .B(n1327), .Z(\mul_a2/fa1_s0[8] ) );
  HS65_GSS_XNOR2X3 U1416 ( .A(n1330), .B(n1329), .Z(\mul_a2/fa1_s0[9] ) );
  HS65_GSS_XNOR2X3 U1417 ( .A(n1332), .B(n1331), .Z(\mul_a2/fa1_s0[10] ) );
  HS65_GSS_XNOR2X3 U1418 ( .A(n1334), .B(n1333), .Z(\mul_a2/fa1_s0[11] ) );
  HS65_GSS_XNOR2X3 U1419 ( .A(n1336), .B(n1335), .Z(\mul_a2/fa1_s0[12] ) );
  HS65_GSS_XNOR2X3 U1420 ( .A(n1338), .B(n1337), .Z(\mul_a2/fa1_s0[13] ) );
  HS65_GSS_XNOR2X3 U1421 ( .A(n1340), .B(n1339), .Z(\mul_a2/fa1_s0[14] ) );
  HS65_GSS_XNOR2X3 U1422 ( .A(n1342), .B(n1341), .Z(\mul_a2/fa1_s0[15] ) );
  HS65_GSS_XNOR2X3 U1423 ( .A(n1344), .B(n1343), .Z(\mul_a2/fa1_s0[16] ) );
  HS65_GS_NOR2X2 U1424 ( .A(y_z2[15]), .B(n1345), .Z(n1347) );
  HS65_GSS_XNOR2X6 U1425 ( .A(n1347), .B(n1346), .Z(\mul_a2/fa1_s0[28] ) );
  HS65_GSS_XNOR2X3 U1426 ( .A(x_z2[15]), .B(n1348), .Z(n1377) );
  HS65_GS_HA1X4 U1427 ( .A0(n1692), .B0(n1349), .CO(n1379), .S0(n1376) );
  HS65_GS_PAO2X4 U1428 ( .A(n1377), .B(n1376), .P(n1712), .Z(
        \mul_b1/fa1_c0[18] ) );
  HS65_GS_HA1X4 U1429 ( .A0(n1680), .B0(n1350), .CO(n1351), .S0(n1627) );
  HS65_GSS_XOR3X2 U1430 ( .A(x_z2[4]), .B(\mul_b1/fa1_s0[0] ), .C(n1627), .Z(
        \mul_b1/fa1_s0[4] ) );
  HS65_GS_HA1X4 U1431 ( .A0(n1679), .B0(n1678), .CO(n1352), .S0(n1629) );
  HS65_GS_HA1X4 U1432 ( .A0(n1681), .B0(n1351), .CO(n1353), .S0(n1628) );
  HS65_GSS_XOR3X2 U1433 ( .A(x_z2[5]), .B(n1629), .C(n1628), .Z(
        \mul_b1/fa1_s0[5] ) );
  HS65_GS_HA1X4 U1434 ( .A0(n1680), .B0(n1352), .CO(n1355), .S0(n1631) );
  HS65_GS_HA1X4 U1435 ( .A0(n1682), .B0(n1353), .CO(n1354), .S0(n1630) );
  HS65_GSS_XOR3X2 U1436 ( .A(x_z2[6]), .B(n1631), .C(n1630), .Z(
        \mul_b1/fa1_s0[6] ) );
  HS65_GS_HA1X4 U1437 ( .A0(n1683), .B0(n1354), .CO(n1356), .S0(n1633) );
  HS65_GS_HA1X4 U1438 ( .A0(n1681), .B0(n1355), .CO(n1357), .S0(n1632) );
  HS65_GSS_XOR3X2 U1439 ( .A(x_z2[7]), .B(n1633), .C(n1632), .Z(
        \mul_b1/fa1_s0[7] ) );
  HS65_GS_HA1X4 U1440 ( .A0(n1684), .B0(n1356), .CO(n1358), .S0(n1635) );
  HS65_GS_HA1X4 U1441 ( .A0(n1682), .B0(n1357), .CO(n1359), .S0(n1634) );
  HS65_GSS_XOR3X2 U1442 ( .A(x_z2[8]), .B(n1635), .C(n1634), .Z(
        \mul_b1/fa1_s0[8] ) );
  HS65_GS_HA1X4 U1443 ( .A0(n1685), .B0(n1358), .CO(n1360), .S0(n1637) );
  HS65_GS_HA1X4 U1444 ( .A0(n1683), .B0(n1359), .CO(n1361), .S0(n1636) );
  HS65_GSS_XOR3X2 U1445 ( .A(x_z2[9]), .B(n1637), .C(n1636), .Z(
        \mul_b1/fa1_s0[9] ) );
  HS65_GS_HA1X4 U1446 ( .A0(n1686), .B0(n1360), .CO(n1362), .S0(n1639) );
  HS65_GS_HA1X4 U1447 ( .A0(n1684), .B0(n1361), .CO(n1363), .S0(n1638) );
  HS65_GSS_XOR3X2 U1448 ( .A(x_z2[10]), .B(n1639), .C(n1638), .Z(
        \mul_b1/fa1_s0[10] ) );
  HS65_GS_HA1X4 U1449 ( .A0(n1687), .B0(n1362), .CO(n1364), .S0(n1641) );
  HS65_GS_HA1X4 U1450 ( .A0(n1685), .B0(n1363), .CO(n1365), .S0(n1640) );
  HS65_GSS_XOR3X2 U1451 ( .A(x_z2[11]), .B(n1641), .C(n1640), .Z(
        \mul_b1/fa1_s0[11] ) );
  HS65_GS_HA1X4 U1452 ( .A0(n1688), .B0(n1364), .CO(n1367), .S0(n1643) );
  HS65_GS_HA1X4 U1453 ( .A0(n1686), .B0(n1365), .CO(n1366), .S0(n1642) );
  HS65_GSS_XOR3X2 U1454 ( .A(x_z2[12]), .B(n1643), .C(n1642), .Z(
        \mul_b1/fa1_s0[12] ) );
  HS65_GS_HA1X4 U1455 ( .A0(n1687), .B0(n1366), .CO(n1368), .S0(n1645) );
  HS65_GS_HA1X4 U1456 ( .A0(n1689), .B0(n1367), .CO(n1369), .S0(n1644) );
  HS65_GSS_XOR3X2 U1457 ( .A(x_z2[13]), .B(n1645), .C(n1644), .Z(
        \mul_b1/fa1_s0[13] ) );
  HS65_GS_HA1X4 U1458 ( .A0(n1688), .B0(n1368), .CO(n1371), .S0(n1647) );
  HS65_GS_HA1X4 U1459 ( .A0(n1690), .B0(n1369), .CO(n1370), .S0(n1646) );
  HS65_GSS_XOR3X2 U1460 ( .A(x_z2[14]), .B(n1647), .C(n1646), .Z(
        \mul_b1/fa1_s0[14] ) );
  HS65_GS_HA1X4 U1461 ( .A0(n1691), .B0(n1370), .CO(n1373), .S0(n1649) );
  HS65_GS_HA1X4 U1462 ( .A0(n1689), .B0(n1371), .CO(n1372), .S0(n1648) );
  HS65_GSS_XOR3X2 U1463 ( .A(x_z2[15]), .B(n1649), .C(n1648), .Z(
        \mul_b1/fa1_s0[15] ) );
  HS65_GS_HA1X4 U1464 ( .A0(n1690), .B0(n1372), .CO(n1375), .S0(n1651) );
  HS65_GS_HA1X4 U1465 ( .A0(n1692), .B0(n1373), .CO(n1374), .S0(n1650) );
  HS65_GSS_XOR3X2 U1466 ( .A(x_z2[15]), .B(n1651), .C(n1650), .Z(
        \mul_b1/fa1_s0[16] ) );
  HS65_GS_HA1X4 U1467 ( .A0(n1693), .B0(n1374), .CO(n1348), .S0(n1408) );
  HS65_GS_HA1X4 U1468 ( .A0(n1691), .B0(n1375), .CO(n1349), .S0(n1407) );
  HS65_GSS_XOR3X2 U1469 ( .A(x_z2[15]), .B(n1408), .C(n1407), .Z(
        \mul_b1/fa1_s0[17] ) );
  HS65_GSS_XOR3X2 U1470 ( .A(x_z2[15]), .B(n1377), .C(n1376), .Z(
        \mul_b1/fa1_s0[18] ) );
  HS65_GSS_XNOR2X3 U1471 ( .A(n2), .B(n1693), .Z(n1383) );
  HS65_GSS_XNOR2X3 U1472 ( .A(n1383), .B(n1378), .Z(\mul_b1/fa1_s0[19] ) );
  HS65_GS_HA1X4 U1473 ( .A0(n1693), .B0(n1379), .CO(n1381), .S0(n930) );
  HS65_GSS_XOR2X3 U1474 ( .A(x_z2[15]), .B(n1381), .Z(n1380) );
  HS65_GSS_XNOR2X3 U1475 ( .A(n1383), .B(n1380), .Z(\mul_b1/fa1_s0[20] ) );
  HS65_GS_OR2X4 U1476 ( .A(x_z2[15]), .B(n1381), .Z(n1382) );
  HS65_GSS_XNOR2X3 U1477 ( .A(n1383), .B(n1382), .Z(\mul_b1/fa1_s0[28] ) );
  HS65_GS_AND2X4 U1478 ( .A(n1610), .B(\mul_b1/fa1_s0[0] ), .Z(
        \mul_b1/fa1_c2[14] ) );
  HS65_GS_HA1X4 U1479 ( .A0(n1679), .B0(n1678), .CO(n1384), .S0(n1610) );
  HS65_GS_AND2X4 U1480 ( .A(n1611), .B(\mul_b1/fa1_s0[1] ), .Z(
        \mul_b1/fa1_c2[15] ) );
  HS65_GS_HA1X4 U1481 ( .A0(n1680), .B0(n1384), .CO(n1385), .S0(n1611) );
  HS65_GS_AND2X4 U1482 ( .A(n1612), .B(x_z2[2]), .Z(\mul_b1/fa1_c2[16] ) );
  HS65_GS_HA1X4 U1483 ( .A0(n1681), .B0(n1385), .CO(n1386), .S0(n1612) );
  HS65_GS_AND2X4 U1484 ( .A(n1613), .B(x_z2[3]), .Z(\mul_b1/fa1_c2[17] ) );
  HS65_GS_HA1X4 U1485 ( .A0(n1682), .B0(n1386), .CO(n1387), .S0(n1613) );
  HS65_GS_AND2X4 U1486 ( .A(n1614), .B(x_z2[4]), .Z(\mul_b1/fa1_c2[18] ) );
  HS65_GS_HA1X4 U1487 ( .A0(n1683), .B0(n1387), .CO(n1388), .S0(n1614) );
  HS65_GS_AND2X4 U1488 ( .A(n1615), .B(x_z2[5]), .Z(\mul_b1/fa1_c2[19] ) );
  HS65_GS_HA1X4 U1489 ( .A0(n1684), .B0(n1388), .CO(n1389), .S0(n1615) );
  HS65_GS_AND2X4 U1490 ( .A(n1616), .B(x_z2[6]), .Z(\mul_b1/fa1_c2[20] ) );
  HS65_GS_HA1X4 U1491 ( .A0(n1685), .B0(n1389), .CO(n1390), .S0(n1616) );
  HS65_GS_AND2X4 U1492 ( .A(n1617), .B(x_z2[7]), .Z(\mul_b1/fa1_c2[21] ) );
  HS65_GS_HA1X4 U1493 ( .A0(n1686), .B0(n1390), .CO(n1391), .S0(n1617) );
  HS65_GS_AND2X4 U1494 ( .A(n1618), .B(x_z2[8]), .Z(\mul_b1/fa1_c2[22] ) );
  HS65_GS_HA1X4 U1495 ( .A0(n1687), .B0(n1391), .CO(n1392), .S0(n1618) );
  HS65_GS_AND2X4 U1496 ( .A(n1619), .B(x_z2[9]), .Z(\mul_b1/fa1_c2[23] ) );
  HS65_GS_HA1X4 U1497 ( .A0(n1688), .B0(n1392), .CO(n1393), .S0(n1619) );
  HS65_GS_AND2X4 U1498 ( .A(n1620), .B(x_z2[10]), .Z(\mul_b1/fa1_c2[24] ) );
  HS65_GS_HA1X4 U1499 ( .A0(n1689), .B0(n1393), .CO(n1394), .S0(n1620) );
  HS65_GS_AND2X4 U1500 ( .A(n1621), .B(x_z2[11]), .Z(\mul_b1/fa1_c2[25] ) );
  HS65_GS_HA1X4 U1501 ( .A0(n1690), .B0(n1394), .CO(n1395), .S0(n1621) );
  HS65_GS_AND2X4 U1502 ( .A(n1622), .B(x_z2[12]), .Z(\mul_b1/fa1_c2[26] ) );
  HS65_GS_HA1X4 U1503 ( .A0(n1691), .B0(n1395), .CO(n1396), .S0(n1622) );
  HS65_GS_AND2X4 U1504 ( .A(n1623), .B(x_z2[13]), .Z(\mul_b1/fa1_c2[27] ) );
  HS65_GS_HA1X4 U1505 ( .A0(n1692), .B0(n1396), .CO(n1625), .S0(n1623) );
  HS65_GSS_XNOR2X3 U1506 ( .A(n1712), .B(n1625), .Z(n1624) );
  HS65_GS_AND2X4 U1507 ( .A(n1624), .B(x_z2[14]), .Z(\mul_b1/fa1_c2[28] ) );
  HS65_GS_AOI12X2 U1508 ( .A(n1400), .B(n1399), .C(n1397), .Z(n1398) );
  HS65_GS_CB4I6X4 U1509 ( .A(n1400), .B(n1399), .C(n1398), .D(n1404), .Z(
        \mul_b2/result_sat[13] ) );
  HS65_GS_FA1X4 U1510 ( .A0(n1403), .B0(n1402), .CI(n1401), .CO(n937), .S0(
        n1406) );
  HS65_GS_AO12X4 U1511 ( .A(n1406), .B(n1405), .C(n1404), .Z(
        \mul_b2/result_sat[14] ) );
  HS65_GS_PAO2X4 U1512 ( .A(n1408), .B(n1407), .P(x_z2[15]), .Z(
        \mul_b1/fa1_c0[17] ) );
  HS65_GS_AOI12X2 U1513 ( .A(n1411), .B(n1410), .C(n1436), .Z(n1409) );
  HS65_GS_CB4I6X4 U1514 ( .A(n1411), .B(n1410), .C(n1409), .D(n1443), .Z(
        \mul_a1/result_sat[1] ) );
  HS65_GS_FA1X4 U1515 ( .A0(n1414), .B0(n1413), .CI(n1412), .CO(n1416), .S0(
        n1415) );
  HS65_GS_AO12X4 U1516 ( .A(n1415), .B(n1444), .C(n1443), .Z(
        \mul_a1/result_sat[2] ) );
  HS65_GS_FA1X4 U1517 ( .A0(n1418), .B0(n1417), .CI(n1416), .CO(n1422), .S0(
        n1419) );
  HS65_GS_AO12X4 U1518 ( .A(n1419), .B(n1444), .C(n1443), .Z(
        \mul_a1/result_sat[3] ) );
  HS65_GS_FA1X4 U1519 ( .A0(n1422), .B0(n1421), .CI(n1420), .CO(n1426), .S0(
        n1423) );
  HS65_GS_AO12X4 U1520 ( .A(n1423), .B(n1444), .C(n1443), .Z(
        \mul_a1/result_sat[4] ) );
  HS65_GS_FA1X4 U1521 ( .A0(n1426), .B0(n1425), .CI(n1424), .CO(n1430), .S0(
        n1427) );
  HS65_GS_AO12X4 U1522 ( .A(n1427), .B(n1444), .C(n1443), .Z(
        \mul_a1/result_sat[5] ) );
  HS65_GS_FA1X4 U1523 ( .A0(n1430), .B0(n1429), .CI(n1428), .CO(n1434), .S0(
        n1431) );
  HS65_GS_AO12X4 U1524 ( .A(n1431), .B(n1444), .C(n1443), .Z(
        \mul_a1/result_sat[6] ) );
  HS65_GS_FA1X4 U1525 ( .A0(n1434), .B0(n1433), .CI(n1432), .CO(n1029), .S0(
        n1435) );
  HS65_GS_AO12X4 U1526 ( .A(n1435), .B(n1444), .C(n1443), .Z(
        \mul_a1/result_sat[7] ) );
  HS65_GS_AOI12X2 U1527 ( .A(n1439), .B(n1438), .C(n1436), .Z(n1437) );
  HS65_GS_CB4I6X4 U1528 ( .A(n1439), .B(n1438), .C(n1437), .D(n1443), .Z(
        \mul_a1/result_sat[13] ) );
  HS65_GS_FA1X4 U1529 ( .A0(n1442), .B0(n1441), .CI(n1440), .CO(n1013), .S0(
        n1445) );
  HS65_GS_AO12X4 U1530 ( .A(n1445), .B(n1444), .C(n1443), .Z(
        \mul_a1/result_sat[14] ) );
  HS65_GS_AND2X4 U1531 ( .A(y_z1[2]), .B(y_z1[0]), .Z(\mul_a1/fa1_c1[8] ) );
  HS65_GS_HA1X4 U1532 ( .A0(n1447), .B0(n1446), .CO(n1448), .S0(n1485) );
  HS65_GS_AND2X4 U1533 ( .A(y_z1[3]), .B(n1485), .Z(\mul_a1/fa1_c1[9] ) );
  HS65_GS_HA1X4 U1534 ( .A0(n1484), .B0(n1448), .CO(n1451), .S0(n1486) );
  HS65_GS_IVX2 U1535 ( .A(n1486), .Z(n1450) );
  HS65_GS_OAI21X2 U1536 ( .A(y_z1[4]), .B(n1486), .C(y_z1[0]), .Z(n1449) );
  HS65_GS_OAI21X2 U1537 ( .A(n1675), .B(n1450), .C(n1449), .Z(
        \mul_a1/fa1_c1[10] ) );
  HS65_GS_HA1X4 U1538 ( .A0(n1677), .B0(n1451), .CO(n1454), .S0(n1487) );
  HS65_GS_IVX2 U1539 ( .A(n1487), .Z(n1453) );
  HS65_GS_OAI21X2 U1540 ( .A(y_z1[5]), .B(n1487), .C(y_z1[1]), .Z(n1452) );
  HS65_GS_OAI21X2 U1541 ( .A(n1673), .B(n1453), .C(n1452), .Z(
        \mul_a1/fa1_c1[11] ) );
  HS65_GS_HA1X4 U1542 ( .A0(n1675), .B0(n1454), .CO(n1457), .S0(n1488) );
  HS65_GS_IVX2 U1543 ( .A(n1488), .Z(n1456) );
  HS65_GS_OAI21X2 U1544 ( .A(y_z1[6]), .B(n1488), .C(y_z1[2]), .Z(n1455) );
  HS65_GS_OAI21X2 U1545 ( .A(n1671), .B(n1456), .C(n1455), .Z(
        \mul_a1/fa1_c1[12] ) );
  HS65_GS_HA1X4 U1546 ( .A0(n1673), .B0(n1457), .CO(n1460), .S0(n1489) );
  HS65_GS_IVX2 U1547 ( .A(n1489), .Z(n1459) );
  HS65_GS_OAI21X2 U1548 ( .A(y_z1[7]), .B(n1489), .C(y_z1[3]), .Z(n1458) );
  HS65_GS_OAI21X2 U1549 ( .A(n1669), .B(n1459), .C(n1458), .Z(
        \mul_a1/fa1_c1[13] ) );
  HS65_GS_HA1X4 U1550 ( .A0(n1671), .B0(n1460), .CO(n1463), .S0(n1490) );
  HS65_GS_IVX2 U1551 ( .A(n1490), .Z(n1462) );
  HS65_GS_OAI21X2 U1552 ( .A(y_z1[8]), .B(n1490), .C(y_z1[4]), .Z(n1461) );
  HS65_GS_OAI21X2 U1553 ( .A(n1667), .B(n1462), .C(n1461), .Z(
        \mul_a1/fa1_c1[14] ) );
  HS65_GS_HA1X4 U1554 ( .A0(n1669), .B0(n1463), .CO(n1466), .S0(n1491) );
  HS65_GS_IVX2 U1555 ( .A(n1491), .Z(n1465) );
  HS65_GS_OAI21X2 U1556 ( .A(y_z1[9]), .B(n1491), .C(y_z1[5]), .Z(n1464) );
  HS65_GS_OAI21X2 U1557 ( .A(n1665), .B(n1465), .C(n1464), .Z(
        \mul_a1/fa1_c1[15] ) );
  HS65_GS_HA1X4 U1558 ( .A0(n1667), .B0(n1466), .CO(n1469), .S0(n1492) );
  HS65_GS_IVX2 U1559 ( .A(n1492), .Z(n1468) );
  HS65_GS_OAI21X2 U1560 ( .A(y_z1[10]), .B(n1492), .C(y_z1[6]), .Z(n1467) );
  HS65_GS_OAI21X2 U1561 ( .A(n1663), .B(n1468), .C(n1467), .Z(
        \mul_a1/fa1_c1[16] ) );
  HS65_GS_HA1X4 U1562 ( .A0(n1665), .B0(n1469), .CO(n1046), .S0(n1493) );
  HS65_GS_IVX2 U1563 ( .A(n1493), .Z(n1471) );
  HS65_GS_OAI21X2 U1564 ( .A(y_z1[11]), .B(n1493), .C(y_z1[7]), .Z(n1470) );
  HS65_GS_OAI21X2 U1565 ( .A(n1661), .B(n1471), .C(n1470), .Z(
        \mul_a1/fa1_c1[17] ) );
  HS65_GS_HA1X4 U1566 ( .A0(n1661), .B0(n1472), .CO(n1049), .S0(n1495) );
  HS65_GS_IVX2 U1567 ( .A(n1495), .Z(n1474) );
  HS65_GS_OAI21X2 U1568 ( .A(y_z1[13]), .B(n1495), .C(y_z1[9]), .Z(n1473) );
  HS65_GS_OAI21X2 U1569 ( .A(n1657), .B(n1474), .C(n1473), .Z(
        \mul_a1/fa1_c1[19] ) );
  HS65_GS_HA1X4 U1570 ( .A0(n1657), .B0(n1475), .CO(n1478), .S0(n1497) );
  HS65_GS_IVX2 U1571 ( .A(n1497), .Z(n1477) );
  HS65_GS_OAI21X2 U1572 ( .A(y_z1[15]), .B(n1497), .C(y_z1[11]), .Z(n1476) );
  HS65_GS_OAI21X2 U1573 ( .A(n1483), .B(n1477), .C(n1476), .Z(
        \mul_a1/fa1_c1[21] ) );
  HS65_GS_HA1X4 U1574 ( .A0(n1655), .B0(n1478), .CO(n1481), .S0(n1498) );
  HS65_GS_IVX2 U1575 ( .A(n1498), .Z(n1480) );
  HS65_GS_OAI21X2 U1576 ( .A(y_z1[15]), .B(n1498), .C(y_z1[12]), .Z(n1479) );
  HS65_GS_OAI21X2 U1577 ( .A(n1483), .B(n1480), .C(n1479), .Z(
        \mul_a1/fa1_c1[22] ) );
  HS65_GS_HA1X4 U1578 ( .A0(n1483), .B0(n1481), .CO(n1500), .S0(n1499) );
  HS65_GS_IVX2 U1579 ( .A(n1499), .Z(n1482) );
  HS65_GS_OAI21X2 U1580 ( .A(n1483), .B(n1482), .C(n1657), .Z(
        \mul_a1/fa1_c1[23] ) );
  HS65_GSS_XNOR2X3 U1581 ( .A(y_z1[0]), .B(n1484), .Z(\mul_a1/fa1_s1[8] ) );
  HS65_GSS_XNOR2X3 U1582 ( .A(n1485), .B(n1677), .Z(\mul_a1/fa1_s1[9] ) );
  HS65_GSS_XOR3X2 U1583 ( .A(y_z1[0]), .B(y_z1[4]), .C(n1486), .Z(
        \mul_a1/fa1_s1[10] ) );
  HS65_GSS_XOR3X2 U1584 ( .A(y_z1[5]), .B(y_z1[1]), .C(n1487), .Z(
        \mul_a1/fa1_s1[11] ) );
  HS65_GSS_XOR3X2 U1585 ( .A(y_z1[6]), .B(y_z1[2]), .C(n1488), .Z(
        \mul_a1/fa1_s1[12] ) );
  HS65_GSS_XOR3X2 U1586 ( .A(y_z1[3]), .B(y_z1[7]), .C(n1489), .Z(
        \mul_a1/fa1_s1[13] ) );
  HS65_GSS_XOR3X2 U1587 ( .A(y_z1[4]), .B(y_z1[8]), .C(n1490), .Z(
        \mul_a1/fa1_s1[14] ) );
  HS65_GSS_XOR3X2 U1588 ( .A(y_z1[5]), .B(y_z1[9]), .C(n1491), .Z(
        \mul_a1/fa1_s1[15] ) );
  HS65_GSS_XOR3X2 U1589 ( .A(y_z1[6]), .B(y_z1[10]), .C(n1492), .Z(
        \mul_a1/fa1_s1[16] ) );
  HS65_GSS_XOR3X2 U1590 ( .A(y_z1[7]), .B(y_z1[11]), .C(n1493), .Z(
        \mul_a1/fa1_s1[17] ) );
  HS65_GSS_XOR3X2 U1591 ( .A(y_z1[8]), .B(y_z1[12]), .C(n1494), .Z(
        \mul_a1/fa1_s1[18] ) );
  HS65_GSS_XOR3X2 U1592 ( .A(y_z1[9]), .B(y_z1[13]), .C(n1495), .Z(
        \mul_a1/fa1_s1[19] ) );
  HS65_GSS_XOR3X2 U1593 ( .A(y_z1[14]), .B(y_z1[10]), .C(n1496), .Z(
        \mul_a1/fa1_s1[20] ) );
  HS65_GSS_XOR3X2 U1594 ( .A(y_z1[15]), .B(y_z1[11]), .C(n1497), .Z(
        \mul_a1/fa1_s1[21] ) );
  HS65_GSS_XOR3X2 U1595 ( .A(y_z1[15]), .B(y_z1[12]), .C(n1498), .Z(
        \mul_a1/fa1_s1[22] ) );
  HS65_GSS_XOR3X2 U1596 ( .A(y_z1[15]), .B(y_z1[13]), .C(n1499), .Z(
        \mul_a1/fa1_s1[23] ) );
  HS65_GSS_XNOR2X3 U1597 ( .A(y_z1[15]), .B(n1500), .Z(n1501) );
  HS65_GSS_XOR3X2 U1598 ( .A(n1501), .B(y_z1[14]), .C(y_z1[15]), .Z(
        \mul_a1/fa1_s1[24] ) );
  HS65_GS_AOI12X2 U1599 ( .A(n1505), .B(n1504), .C(n1502), .Z(n1503) );
  HS65_GS_CB4I6X4 U1600 ( .A(n1505), .B(n1504), .C(n1503), .D(n1509), .Z(
        \mul_b0/result_sat[13] ) );
  HS65_GS_FA1X4 U1601 ( .A0(n1508), .B0(n1507), .CI(n1506), .CO(n1063), .S0(
        n1511) );
  HS65_GS_AO12X4 U1602 ( .A(n1511), .B(n1510), .C(n1509), .Z(
        \mul_b0/result_sat[14] ) );
  HS65_GS_AND2X4 U1603 ( .A(x_z1[5]), .B(x_z1[0]), .Z(\mul_b0/fa1_c0[5] ) );
  HS65_GS_HA1X4 U1604 ( .A0(n1513), .B0(n1512), .CO(n1514), .S0(n1533) );
  HS65_GS_AND2X4 U1605 ( .A(n1533), .B(x_z1[6]), .Z(\mul_b0/fa1_c0[6] ) );
  HS65_GS_HA1X4 U1606 ( .A0(n1515), .B0(n1514), .CO(n1516), .S0(n1535) );
  HS65_GS_AND2X4 U1607 ( .A(x_z1[7]), .B(n1535), .Z(\mul_b0/fa1_c0[7] ) );
  HS65_GS_HA1X4 U1608 ( .A0(n1517), .B0(n1516), .CO(n1518), .S0(n1537) );
  HS65_GS_AND2X4 U1609 ( .A(n1537), .B(x_z1[8]), .Z(\mul_b0/fa1_c0[8] ) );
  HS65_GS_HA1X4 U1610 ( .A0(n1519), .B0(n1518), .CO(n1520), .S0(n1539) );
  HS65_GS_AND2X4 U1611 ( .A(n1539), .B(x_z1[9]), .Z(\mul_b0/fa1_c0[9] ) );
  HS65_GS_HA1X4 U1612 ( .A0(n1521), .B0(n1520), .CO(n1522), .S0(n1541) );
  HS65_GS_AND2X4 U1613 ( .A(n1541), .B(x_z1[10]), .Z(\mul_b0/fa1_c0[10] ) );
  HS65_GS_HA1X4 U1614 ( .A0(n1532), .B0(n1522), .CO(n1523), .S0(n1543) );
  HS65_GS_AND2X4 U1615 ( .A(n1543), .B(x_z1[11]), .Z(\mul_b0/fa1_c0[11] ) );
  HS65_GS_HA1X4 U1616 ( .A0(n1534), .B0(n1523), .CO(n1524), .S0(n1545) );
  HS65_GS_AND2X4 U1617 ( .A(n1545), .B(x_z1[12]), .Z(\mul_b0/fa1_c0[12] ) );
  HS65_GS_HA1X4 U1618 ( .A0(n1536), .B0(n1524), .CO(n1525), .S0(n1547) );
  HS65_GS_AND2X4 U1619 ( .A(n1547), .B(x_z1[13]), .Z(\mul_b0/fa1_c0[13] ) );
  HS65_GS_HA1X4 U1620 ( .A0(n1538), .B0(n1525), .CO(n1526), .S0(n1549) );
  HS65_GS_AND2X4 U1621 ( .A(n1549), .B(x_z1[14]), .Z(\mul_b0/fa1_c0[14] ) );
  HS65_GS_HA1X4 U1622 ( .A0(n1540), .B0(n1526), .CO(n1527), .S0(n1550) );
  HS65_GS_AND2X4 U1623 ( .A(n1550), .B(n1713), .Z(\mul_b0/fa1_c0[15] ) );
  HS65_GS_HA1X4 U1624 ( .A0(n1542), .B0(n1527), .CO(n1528), .S0(n1551) );
  HS65_GS_AND2X4 U1625 ( .A(n1551), .B(x_z1[15]), .Z(\mul_b0/fa1_c0[16] ) );
  HS65_GS_HA1X4 U1626 ( .A0(n1544), .B0(n1528), .CO(n1529), .S0(n1552) );
  HS65_GS_AND2X4 U1627 ( .A(n1552), .B(n1713), .Z(\mul_b0/fa1_c0[17] ) );
  HS65_GS_HA1X4 U1628 ( .A0(n1546), .B0(n1529), .CO(n1530), .S0(n1553) );
  HS65_GS_AND2X4 U1629 ( .A(n1553), .B(x_z1[15]), .Z(\mul_b0/fa1_c0[18] ) );
  HS65_GS_HA1X4 U1630 ( .A0(n1548), .B0(n1530), .CO(n1154), .S0(n1555) );
  HS65_GS_AND2X4 U1631 ( .A(n1555), .B(n1713), .Z(\mul_b0/fa1_c0[19] ) );
  HS65_GS_AND2X4 U1632 ( .A(n1531), .B(x_z1[15]), .Z(\mul_b0/fa1_c0[20] ) );
  HS65_GSS_XNOR2X3 U1633 ( .A(n1533), .B(n1532), .Z(\mul_b0/fa1_s0[6] ) );
  HS65_GSS_XNOR2X3 U1634 ( .A(n1535), .B(n1534), .Z(\mul_b0/fa1_s0[7] ) );
  HS65_GSS_XNOR2X3 U1635 ( .A(n1537), .B(n1536), .Z(\mul_b0/fa1_s0[8] ) );
  HS65_GSS_XNOR2X3 U1636 ( .A(n1539), .B(n1538), .Z(\mul_b0/fa1_s0[9] ) );
  HS65_GSS_XNOR2X3 U1637 ( .A(n1541), .B(n1540), .Z(\mul_b0/fa1_s0[10] ) );
  HS65_GSS_XNOR2X3 U1638 ( .A(n1543), .B(n1542), .Z(\mul_b0/fa1_s0[11] ) );
  HS65_GSS_XNOR2X3 U1639 ( .A(n1545), .B(n1544), .Z(\mul_b0/fa1_s0[12] ) );
  HS65_GSS_XNOR2X3 U1640 ( .A(n1547), .B(n1546), .Z(\mul_b0/fa1_s0[13] ) );
  HS65_GSS_XNOR2X3 U1641 ( .A(n1549), .B(n1548), .Z(\mul_b0/fa1_s0[14] ) );
  HS65_GSS_XNOR2X3 U1642 ( .A(n1550), .B(n1554), .Z(\mul_b0/fa1_s0[15] ) );
  HS65_GSS_XNOR2X3 U1643 ( .A(n1551), .B(n1554), .Z(\mul_b0/fa1_s0[16] ) );
  HS65_GSS_XNOR2X3 U1644 ( .A(n1552), .B(n1554), .Z(\mul_b0/fa1_s0[17] ) );
  HS65_GSS_XNOR2X3 U1645 ( .A(n1553), .B(n1554), .Z(\mul_b0/fa1_s0[18] ) );
  HS65_GSS_XNOR2X3 U1646 ( .A(n1555), .B(n1554), .Z(\mul_b0/fa1_s0[19] ) );
  HS65_GS_FA1X4 U1647 ( .A0(n1558), .B0(n1557), .CI(n1556), .CO(n1561), .S0(
        n1559) );
  HS65_GS_AO12X4 U1648 ( .A(n1559), .B(n1607), .C(n1609), .Z(
        \mul_b1/result_sat[1] ) );
  HS65_GS_FA1X4 U1649 ( .A0(n1562), .B0(n1561), .CI(n1560), .CO(n1566), .S0(
        n1563) );
  HS65_GS_AO12X4 U1650 ( .A(n1563), .B(n1607), .C(n1609), .Z(
        \mul_b1/result_sat[2] ) );
  HS65_GS_FA1X4 U1651 ( .A0(n1566), .B0(n1565), .CI(n1564), .CO(n1570), .S0(
        n1567) );
  HS65_GS_AO12X4 U1652 ( .A(n1567), .B(n1607), .C(n1609), .Z(
        \mul_b1/result_sat[3] ) );
  HS65_GS_FA1X4 U1653 ( .A0(n1570), .B0(n1569), .CI(n1568), .CO(n1573), .S0(
        n1571) );
  HS65_GS_OA12X4 U1654 ( .A(n1609), .B(n1571), .C(n1607), .Z(
        \mul_b1/result_sat[4] ) );
  HS65_GS_FA1X4 U1655 ( .A0(n1574), .B0(n1573), .CI(n1572), .CO(n1578), .S0(
        n1575) );
  HS65_GS_AO12X4 U1656 ( .A(n1575), .B(n1607), .C(n1609), .Z(
        \mul_b1/result_sat[5] ) );
  HS65_GS_FA1X4 U1657 ( .A0(n1578), .B0(n1577), .CI(n1576), .CO(n1148), .S0(
        n1579) );
  HS65_GS_AO12X4 U1658 ( .A(n1579), .B(n1607), .C(n1609), .Z(
        \mul_b1/result_sat[6] ) );
  HS65_GS_FA1X4 U1659 ( .A0(n1582), .B0(n1581), .CI(n1580), .CO(n1585), .S0(
        n1583) );
  HS65_GS_OA12X4 U1660 ( .A(n1609), .B(n1583), .C(n1607), .Z(
        \mul_b1/result_sat[8] ) );
  HS65_GS_FA1X4 U1661 ( .A0(n1586), .B0(n1585), .CI(n1584), .CO(n1590), .S0(
        n1587) );
  HS65_GS_OA12X4 U1662 ( .A(n1609), .B(n1587), .C(n1607), .Z(
        \mul_b1/result_sat[9] ) );
  HS65_GS_FA1X4 U1663 ( .A0(n1590), .B0(n1589), .CI(n1588), .CO(n1593), .S0(
        n1591) );
  HS65_GS_OA12X4 U1664 ( .A(n1609), .B(n1591), .C(n1607), .Z(
        \mul_b1/result_sat[10] ) );
  HS65_GS_FA1X4 U1665 ( .A0(n1594), .B0(n1593), .CI(n1592), .CO(n1598), .S0(
        n1595) );
  HS65_GS_AO12X4 U1666 ( .A(n1595), .B(n1607), .C(n1609), .Z(
        \mul_b1/result_sat[11] ) );
  HS65_GS_FA1X4 U1667 ( .A0(n1598), .B0(n1597), .CI(n1596), .CO(n1601), .S0(
        n1599) );
  HS65_GS_AO12X4 U1668 ( .A(n1599), .B(n1607), .C(n1609), .Z(
        \mul_b1/result_sat[12] ) );
  HS65_GS_FA1X4 U1669 ( .A0(n1602), .B0(n1601), .CI(n1600), .CO(n1606), .S0(
        n1603) );
  HS65_GS_AO12X4 U1670 ( .A(n1603), .B(n1607), .C(n1609), .Z(
        \mul_b1/result_sat[13] ) );
  HS65_GS_FA1X4 U1671 ( .A0(n1606), .B0(n1605), .CI(n1604), .CO(n1133), .S0(
        n1608) );
  HS65_GS_OA12X4 U1672 ( .A(n1609), .B(n1608), .C(n1607), .Z(
        \mul_b1/result_sat[14] ) );
  HS65_GSS_XNOR2X3 U1673 ( .A(n1610), .B(n1678), .Z(\mul_b1/fa1_s2[14] ) );
  HS65_GSS_XNOR2X3 U1674 ( .A(n1611), .B(n1679), .Z(\mul_b1/fa1_s2[15] ) );
  HS65_GSS_XNOR2X3 U1675 ( .A(n1612), .B(n1680), .Z(\mul_b1/fa1_s2[16] ) );
  HS65_GSS_XNOR2X3 U1676 ( .A(n1613), .B(n1681), .Z(\mul_b1/fa1_s2[17] ) );
  HS65_GSS_XNOR2X3 U1677 ( .A(n1614), .B(n1682), .Z(\mul_b1/fa1_s2[18] ) );
  HS65_GSS_XNOR2X3 U1678 ( .A(n1615), .B(n1683), .Z(\mul_b1/fa1_s2[19] ) );
  HS65_GSS_XNOR2X3 U1679 ( .A(n1616), .B(n1684), .Z(\mul_b1/fa1_s2[20] ) );
  HS65_GSS_XNOR2X3 U1680 ( .A(n1617), .B(n1685), .Z(\mul_b1/fa1_s2[21] ) );
  HS65_GSS_XNOR2X3 U1681 ( .A(n1618), .B(n1686), .Z(\mul_b1/fa1_s2[22] ) );
  HS65_GSS_XNOR2X3 U1682 ( .A(n1619), .B(n1687), .Z(\mul_b1/fa1_s2[23] ) );
  HS65_GSS_XNOR2X3 U1683 ( .A(n1620), .B(n1688), .Z(\mul_b1/fa1_s2[24] ) );
  HS65_GSS_XNOR2X3 U1684 ( .A(n1621), .B(n1689), .Z(\mul_b1/fa1_s2[25] ) );
  HS65_GSS_XNOR2X3 U1685 ( .A(n1622), .B(n1690), .Z(\mul_b1/fa1_s2[26] ) );
  HS65_GSS_XNOR2X3 U1686 ( .A(n1623), .B(n1691), .Z(\mul_b1/fa1_s2[27] ) );
  HS65_GSS_XNOR2X3 U1687 ( .A(n1624), .B(n1692), .Z(\mul_b1/fa1_s2[28] ) );
  HS65_GS_NOR2X2 U1688 ( .A(x_z2[15]), .B(n1625), .Z(n1626) );
  HS65_GSS_XNOR2X3 U1689 ( .A(n1626), .B(n1693), .Z(\mul_b1/fa1_s2[29] ) );
  HS65_GS_PAO2X4 U1690 ( .A(\mul_b1/fa1_s0[0] ), .B(n1627), .P(x_z2[4]), .Z(
        \mul_b1/fa1_c0[4] ) );
  HS65_GS_PAO2X4 U1691 ( .A(n1629), .B(n1628), .P(x_z2[5]), .Z(
        \mul_b1/fa1_c0[5] ) );
  HS65_GS_PAO2X4 U1692 ( .A(n1631), .B(n1630), .P(x_z2[6]), .Z(
        \mul_b1/fa1_c0[6] ) );
  HS65_GS_PAO2X4 U1693 ( .A(n1633), .B(n1632), .P(x_z2[7]), .Z(
        \mul_b1/fa1_c0[7] ) );
  HS65_GS_PAO2X4 U1694 ( .A(n1635), .B(n1634), .P(x_z2[8]), .Z(
        \mul_b1/fa1_c0[8] ) );
  HS65_GS_PAO2X4 U1695 ( .A(n1637), .B(n1636), .P(x_z2[9]), .Z(
        \mul_b1/fa1_c0[9] ) );
  HS65_GS_PAO2X4 U1696 ( .A(n1639), .B(n1638), .P(x_z2[10]), .Z(
        \mul_b1/fa1_c0[10] ) );
  HS65_GS_PAO2X4 U1697 ( .A(n1641), .B(n1640), .P(x_z2[11]), .Z(
        \mul_b1/fa1_c0[11] ) );
  HS65_GS_PAO2X4 U1698 ( .A(n1643), .B(n1642), .P(x_z2[12]), .Z(
        \mul_b1/fa1_c0[12] ) );
  HS65_GS_PAO2X4 U1699 ( .A(n1645), .B(n1644), .P(x_z2[13]), .Z(
        \mul_b1/fa1_c0[13] ) );
  HS65_GS_PAO2X4 U1700 ( .A(n1647), .B(n1646), .P(x_z2[14]), .Z(
        \mul_b1/fa1_c0[14] ) );
  HS65_GS_PAO2X4 U1701 ( .A(n1649), .B(n1648), .P(n1712), .Z(
        \mul_b1/fa1_c0[15] ) );
  HS65_GS_PAO2X4 U1702 ( .A(n1651), .B(n1650), .P(x_z2[15]), .Z(
        \mul_b1/fa1_c0[16] ) );
  HS65_GS_AND2X4 U1703 ( .A(x_z2[3]), .B(n1652), .Z(n1709) );
  HS65_GS_AND2X4 U1704 ( .A(x_z2[2]), .B(\mul_b1/fa1_s0[0] ), .Z(n1710) );
  HS65_GSS_XNOR2X3 U1705 ( .A(y_z1[15]), .B(n1653), .Z(\C50/DATA4_18 ) );
  HS65_GS_HA1X4 U1706 ( .A0(n1655), .B0(n1654), .CO(n1653), .S0(\C50/DATA4_17 ) );
  HS65_GS_HA1X4 U1707 ( .A0(n1657), .B0(n1656), .CO(n1654), .S0(\C50/DATA4_16 ) );
  HS65_GS_HA1X4 U1708 ( .A0(n1659), .B0(n1658), .CO(n1656), .S0(\C50/DATA4_15 ) );
  HS65_GS_HA1X4 U1709 ( .A0(n1661), .B0(n1660), .CO(n1658), .S0(\C50/DATA4_14 ) );
  HS65_GS_HA1X4 U1710 ( .A0(n1663), .B0(n1662), .CO(n1660), .S0(\C50/DATA4_13 ) );
  HS65_GS_HA1X4 U1711 ( .A0(n1665), .B0(n1664), .CO(n1662), .S0(\C50/DATA4_12 ) );
  HS65_GS_HA1X4 U1712 ( .A0(n1667), .B0(n1666), .CO(n1664), .S0(\C50/DATA4_11 ) );
  HS65_GS_HA1X4 U1713 ( .A0(n1669), .B0(n1668), .CO(n1666), .S0(\C50/DATA4_10 ) );
  HS65_GS_HA1X4 U1714 ( .A0(n1671), .B0(n1670), .CO(n1668), .S0(\C50/DATA4_9 )
         );
  HS65_GS_HA1X4 U1715 ( .A0(n1673), .B0(n1672), .CO(n1670), .S0(\C50/DATA4_8 )
         );
  HS65_GS_HA1X4 U1716 ( .A0(n1675), .B0(n1674), .CO(n1672), .S0(\C50/DATA4_7 )
         );
  HS65_GS_HA1X4 U1717 ( .A0(n1677), .B0(n1676), .CO(n1674), .S0(\C50/DATA4_6 )
         );
  HS65_GS_AOI12X2 U1718 ( .A(n1678), .B(n1680), .C(\mul_b1/fa1_c1[8] ), .Z(
        \mul_b1/fa1_s1[8] ) );
  HS65_GS_AOI12X2 U1719 ( .A(n1679), .B(n1681), .C(\mul_b1/fa1_c1[9] ), .Z(
        \mul_b1/fa1_s1[9] ) );
  HS65_GS_AOI12X2 U1720 ( .A(n1680), .B(n1682), .C(\mul_b1/fa1_c1[10] ), .Z(
        \mul_b1/fa1_s1[10] ) );
  HS65_GS_AOI12X2 U1721 ( .A(n1681), .B(n1683), .C(\mul_b1/fa1_c1[11] ), .Z(
        \mul_b1/fa1_s1[11] ) );
  HS65_GS_AOI12X2 U1722 ( .A(n1682), .B(n1684), .C(\mul_b1/fa1_c1[12] ), .Z(
        \mul_b1/fa1_s1[12] ) );
  HS65_GS_AOI12X2 U1723 ( .A(n1683), .B(n1685), .C(\mul_b1/fa1_c1[13] ), .Z(
        \mul_b1/fa1_s1[13] ) );
  HS65_GS_AOI12X2 U1724 ( .A(n1684), .B(n1686), .C(\mul_b1/fa1_c1[14] ), .Z(
        \mul_b1/fa1_s1[14] ) );
  HS65_GS_AOI12X2 U1725 ( .A(n1685), .B(n1687), .C(\mul_b1/fa1_c1[15] ), .Z(
        \mul_b1/fa1_s1[15] ) );
  HS65_GS_AOI12X2 U1726 ( .A(n1686), .B(n1688), .C(\mul_b1/fa1_c1[16] ), .Z(
        \mul_b1/fa1_s1[16] ) );
  HS65_GS_AOI12X2 U1727 ( .A(n1687), .B(n1689), .C(\mul_b1/fa1_c1[17] ), .Z(
        \mul_b1/fa1_s1[17] ) );
  HS65_GS_AOI12X2 U1728 ( .A(n1688), .B(n1690), .C(\mul_b1/fa1_c1[18] ), .Z(
        \mul_b1/fa1_s1[18] ) );
  HS65_GS_AOI12X2 U1729 ( .A(n1689), .B(n1691), .C(\mul_b1/fa1_c1[19] ), .Z(
        \mul_b1/fa1_s1[19] ) );
  HS65_GS_AOI12X2 U1730 ( .A(n1690), .B(n1692), .C(\mul_b1/fa1_c1[20] ), .Z(
        \mul_b1/fa1_s1[20] ) );
  HS65_GS_AOI12X2 U1731 ( .A(n1693), .B(n1691), .C(\mul_b1/fa1_c1[21] ), .Z(
        \mul_b1/fa1_s1[21] ) );
  HS65_GS_AOI12X2 U1732 ( .A(n1693), .B(n1692), .C(\mul_b1/fa1_c1[22] ), .Z(
        \mul_b1/fa1_s1[22] ) );
  HS65_GS_FA1X4 U1733 ( .A0(n1696), .B0(n1695), .CI(n1694), .CO(n1700), .S0(
        n1697) );
  HS65_GS_AOI12X2 U1734 ( .A(n1697), .B(n1702), .C(n1701), .Z(
        \mul_a2/result_sat[13] ) );
  HS65_GS_FA1X4 U1735 ( .A0(n1700), .B0(n1699), .CI(n1698), .CO(n879), .S0(
        n1703) );
  HS65_GS_AOI12X2 U1736 ( .A(n1703), .B(n1702), .C(n1701), .Z(
        \mul_a2/result_sat[14] ) );
  HS65_GS_AOI12X2 U1737 ( .A(n1706), .B(n1705), .C(n1704), .Z(n1763) );
endmodule


module opti_sos_0 ( clk, rst_n, data_in, valid_in, b0, b1, b2, a1, a2, 
        data_out, valid_out );
  input [15:0] data_in;
  input [15:0] b0;
  input [15:0] b1;
  input [15:0] b2;
  input [15:0] a1;
  input [15:0] a2;
  output [15:0] data_out;
  input clk, rst_n, valid_in;
  output valid_out;
  wire   valid_T1, valid_T3, valid_T2, \mul_b0/result_sat[15] ,
         \mul_b0/result_sat[14] , \mul_b0/result_sat[13] ,
         \mul_b0/result_sat[12] , \mul_b0/result_sat[11] ,
         \mul_b0/result_sat[10] , \mul_b0/result_sat[9] ,
         \mul_b0/result_sat[8] , \mul_b0/result_sat[7] ,
         \mul_b0/result_sat[6] , \mul_b0/result_sat[5] ,
         \mul_b0/result_sat[4] , \mul_b0/result_sat[3] ,
         \mul_b0/result_sat[2] , \mul_b0/result_sat[1] ,
         \mul_b0/result_sat[0] , \mul_b0/fa1_s2_r[33] , \mul_b0/fa1_s2_r[32] ,
         \mul_b0/fa1_s2_r[31] , \mul_b0/fa1_s2_r[30] , \mul_b0/fa1_s2_r[29] ,
         \mul_b0/fa1_s2_r[28] , \mul_b0/fa1_s2_r[27] , \mul_b0/fa1_s2_r[26] ,
         \mul_b0/fa1_s2_r[25] , \mul_b0/fa1_s2_r[24] , \mul_b0/fa1_s2_r[23] ,
         \mul_b0/fa1_s2_r[22] , \mul_b0/fa1_s2_r[21] , \mul_b0/fa1_s2_r[20] ,
         \mul_b0/fa1_s2_r[19] , \mul_b0/fa1_s2_r[18] , \mul_b0/fa1_s2_r[17] ,
         \mul_b0/fa1_s2_r[16] , \mul_b0/fa1_s2_r[15] , \mul_b0/fa1_s2_r[14] ,
         \mul_b0/fa1_s2_r[13] , \mul_b0/fa1_s2_r[12] , \mul_b0/fa1_s1_r[33] ,
         \mul_b0/fa1_s1_r[32] , \mul_b0/fa1_s1_r[31] , \mul_b0/fa1_s1_r[30] ,
         \mul_b0/fa1_s1_r[29] , \mul_b0/fa1_s1_r[28] , \mul_b0/fa1_s1_r[27] ,
         \mul_b0/fa1_s1_r[26] , \mul_b0/fa1_s1_r[25] , \mul_b0/fa1_s1_r[24] ,
         \mul_b0/fa1_s1_r[23] , \mul_b0/fa1_s1_r[22] , \mul_b0/fa1_s1_r[21] ,
         \mul_b0/fa1_s1_r[20] , \mul_b0/fa1_s1_r[19] , \mul_b0/fa1_s1_r[18] ,
         \mul_b0/fa1_s1_r[17] , \mul_b0/fa1_s1_r[16] , \mul_b0/fa1_s1_r[15] ,
         \mul_b0/fa1_s1_r[14] , \mul_b0/fa1_s1_r[13] , \mul_b0/fa1_s1_r[12] ,
         \mul_b0/fa1_s1_r[11] , \mul_b0/fa1_s1_r[10] , \mul_b0/fa1_s1_r[9] ,
         \mul_b0/fa1_s1_r[8] , \mul_b0/fa1_c0_r[20] , \mul_b0/fa1_c0_r[19] ,
         \mul_b0/fa1_c0_r[18] , \mul_b0/fa1_c0_r[17] , \mul_b0/fa1_c0_r[16] ,
         \mul_b0/fa1_c0_r[15] , \mul_b0/fa1_c0_r[14] , \mul_b0/fa1_c0_r[13] ,
         \mul_b0/fa1_c0_r[12] , \mul_b0/fa1_c0_r[11] , \mul_b0/fa1_c0_r[10] ,
         \mul_b0/fa1_c0_r[9] , \mul_b0/fa1_c0_r[8] , \mul_b0/fa1_c0_r[7] ,
         \mul_b0/fa1_c0_r[6] , \mul_b0/fa1_c0_r[5] , \mul_b0/fa1_s0_r[33] ,
         \mul_b0/fa1_s0_r[32] , \mul_b0/fa1_s0_r[31] , \mul_b0/fa1_s0_r[30] ,
         \mul_b0/fa1_s0_r[29] , \mul_b0/fa1_s0_r[28] , \mul_b0/fa1_s0_r[27] ,
         \mul_b0/fa1_s0_r[26] , \mul_b0/fa1_s0_r[25] , \mul_b0/fa1_s0_r[24] ,
         \mul_b0/fa1_s0_r[23] , \mul_b0/fa1_s0_r[22] , \mul_b0/fa1_s0_r[21] ,
         \mul_b0/fa1_s0_r[20] , \mul_b0/fa1_s0_r[19] , \mul_b0/fa1_s0_r[18] ,
         \mul_b0/fa1_s0_r[17] , \mul_b0/fa1_s0_r[16] , \mul_b0/fa1_s0_r[15] ,
         \mul_b0/fa1_s0_r[14] , \mul_b0/fa1_s0_r[13] , \mul_b0/fa1_s0_r[12] ,
         \mul_b0/fa1_s0_r[11] , \mul_b0/fa1_s0_r[10] , \mul_b0/fa1_s0_r[9] ,
         \mul_b0/fa1_s0_r[8] , \mul_b0/fa1_s0_r[7] , \mul_b0/fa1_s0_r[6] ,
         \mul_b0/fa1_c0[20] , \mul_b0/fa1_c0[19] , \mul_b0/fa1_c0[18] ,
         \mul_b0/fa1_c0[17] , \mul_b0/fa1_c0[16] , \mul_b0/fa1_c0[15] ,
         \mul_b0/fa1_c0[14] , \mul_b0/fa1_c0[13] , \mul_b0/fa1_c0[12] ,
         \mul_b0/fa1_c0[11] , \mul_b0/fa1_c0[10] , \mul_b0/fa1_c0[9] ,
         \mul_b0/fa1_c0[8] , \mul_b0/fa1_c0[7] , \mul_b0/fa1_c0[6] ,
         \mul_b0/fa1_c0[5] , \mul_b0/fa1_s0[30] , \mul_b0/fa1_s0[20] ,
         \mul_b0/fa1_s0[19] , \mul_b0/fa1_s0[18] , \mul_b0/fa1_s0[17] ,
         \mul_b0/fa1_s0[16] , \mul_b0/fa1_s0[15] , \mul_b0/fa1_s0[14] ,
         \mul_b0/fa1_s0[13] , \mul_b0/fa1_s0[12] , \mul_b0/fa1_s0[11] ,
         \mul_b0/fa1_s0[10] , \mul_b0/fa1_s0[9] , \mul_b0/fa1_s0[8] ,
         \mul_b0/fa1_s0[7] , \mul_b0/fa1_s0[6] , \mul_b1/result_sat[15] ,
         \mul_b1/result_sat[14] , \mul_b1/result_sat[13] ,
         \mul_b1/result_sat[12] , \mul_b1/result_sat[11] ,
         \mul_b1/result_sat[10] , \mul_b1/result_sat[9] ,
         \mul_b1/result_sat[8] , \mul_b1/result_sat[7] ,
         \mul_b1/result_sat[6] , \mul_b1/result_sat[5] ,
         \mul_b1/result_sat[4] , \mul_b1/result_sat[3] ,
         \mul_b1/result_sat[2] , \mul_b1/result_sat[1] ,
         \mul_b1/result_sat[0] , \mul_b1/fa1_s2_r[33] , \mul_b1/fa1_s2_r[32] ,
         \mul_b1/fa1_s2_r[31] , \mul_b1/fa1_s2_r[30] , \mul_b1/fa1_s2_r[29] ,
         \mul_b1/fa1_s2_r[28] , \mul_b1/fa1_s2_r[27] , \mul_b1/fa1_s2_r[26] ,
         \mul_b1/fa1_s2_r[25] , \mul_b1/fa1_s2_r[24] , \mul_b1/fa1_s2_r[23] ,
         \mul_b1/fa1_s2_r[22] , \mul_b1/fa1_s2_r[21] , \mul_b1/fa1_s2_r[20] ,
         \mul_b1/fa1_s2_r[19] , \mul_b1/fa1_s2_r[18] , \mul_b1/fa1_s2_r[17] ,
         \mul_b1/fa1_s2_r[16] , \mul_b1/fa1_s2_r[15] , \mul_b1/fa1_s2_r[14] ,
         \mul_b1/fa1_s2_r[13] , \mul_b1/fa1_s2_r[12] , \mul_b1/fa1_c1_r[32] ,
         \mul_b1/fa1_c1_r[31] , \mul_b1/fa1_c1_r[30] , \mul_b1/fa1_c1_r[29] ,
         \mul_b1/fa1_c1_r[28] , \mul_b1/fa1_c1_r[27] , \mul_b1/fa1_c1_r[26] ,
         \mul_b1/fa1_c1_r[25] , \mul_b1/fa1_c1_r[24] , \mul_b1/fa1_c1_r[23] ,
         \mul_b1/fa1_c1_r[22] , \mul_b1/fa1_c1_r[21] , \mul_b1/fa1_c1_r[20] ,
         \mul_b1/fa1_c1_r[19] , \mul_b1/fa1_c1_r[18] , \mul_b1/fa1_c1_r[17] ,
         \mul_b1/fa1_c1_r[16] , \mul_b1/fa1_c1_r[15] , \mul_b1/fa1_c1_r[14] ,
         \mul_b1/fa1_c1_r[13] , \mul_b1/fa1_c1_r[12] , \mul_b1/fa1_c1_r[11] ,
         \mul_b1/fa1_c1_r[10] , \mul_b1/fa1_c1_r[9] , \mul_b1/fa1_c1_r[8] ,
         \mul_b1/fa1_s1_r[22] , \mul_b1/fa1_s1_r[21] , \mul_b1/fa1_s1_r[20] ,
         \mul_b1/fa1_s1_r[19] , \mul_b1/fa1_s1_r[18] , \mul_b1/fa1_s1_r[17] ,
         \mul_b1/fa1_s1_r[16] , \mul_b1/fa1_s1_r[15] , \mul_b1/fa1_s1_r[14] ,
         \mul_b1/fa1_s1_r[13] , \mul_b1/fa1_s1_r[12] , \mul_b1/fa1_s1_r[11] ,
         \mul_b1/fa1_s1_r[10] , \mul_b1/fa1_s1_r[9] , \mul_b1/fa1_s1_r[8] ,
         \mul_b1/fa1_s1_r[7] , \mul_b1/fa1_c0_r[32] , \mul_b1/fa1_c0_r[31] ,
         \mul_b1/fa1_c0_r[30] , \mul_b1/fa1_c0_r[29] , \mul_b1/fa1_c0_r[28] ,
         \mul_b1/fa1_c0_r[27] , \mul_b1/fa1_c0_r[26] , \mul_b1/fa1_c0_r[25] ,
         \mul_b1/fa1_c0_r[24] , \mul_b1/fa1_c0_r[23] , \mul_b1/fa1_c0_r[22] ,
         \mul_b1/fa1_c0_r[21] , \mul_b1/fa1_c0_r[20] , \mul_b1/fa1_c0_r[19] ,
         \mul_b1/fa1_c0_r[18] , \mul_b1/fa1_c0_r[17] , \mul_b1/fa1_c0_r[16] ,
         \mul_b1/fa1_c0_r[15] , \mul_b1/fa1_c0_r[14] , \mul_b1/fa1_c0_r[13] ,
         \mul_b1/fa1_c0_r[12] , \mul_b1/fa1_c0_r[11] , \mul_b1/fa1_c0_r[10] ,
         \mul_b1/fa1_c0_r[9] , \mul_b1/fa1_c0_r[8] , \mul_b1/fa1_c0_r[7] ,
         \mul_b1/fa1_c0_r[6] , \mul_b1/fa1_c0_r[5] , \mul_b1/fa1_c0_r[4] ,
         \mul_b1/fa1_c0_r[3] , \mul_b1/fa1_s0_r[33] , \mul_b1/fa1_s0_r[32] ,
         \mul_b1/fa1_s0_r[31] , \mul_b1/fa1_s0_r[30] , \mul_b1/fa1_s0_r[29] ,
         \mul_b1/fa1_s0_r[28] , \mul_b1/fa1_s0_r[27] , \mul_b1/fa1_s0_r[26] ,
         \mul_b1/fa1_s0_r[25] , \mul_b1/fa1_s0_r[24] , \mul_b1/fa1_s0_r[23] ,
         \mul_b1/fa1_s0_r[22] , \mul_b1/fa1_s0_r[21] , \mul_b1/fa1_s0_r[20] ,
         \mul_b1/fa1_s0_r[19] , \mul_b1/fa1_s0_r[18] , \mul_b1/fa1_s0_r[17] ,
         \mul_b1/fa1_s0_r[16] , \mul_b1/fa1_s0_r[15] , \mul_b1/fa1_s0_r[14] ,
         \mul_b1/fa1_s0_r[13] , \mul_b1/fa1_s0_r[12] , \mul_b1/fa1_s0_r[11] ,
         \mul_b1/fa1_s0_r[10] , \mul_b1/fa1_s0_r[9] , \mul_b1/fa1_s0_r[8] ,
         \mul_b1/fa1_s0_r[7] , \mul_b1/fa1_s0_r[6] , \mul_b1/fa1_s0_r[5] ,
         \mul_b1/fa1_s0_r[4] , \mul_b1/fa1_c1[22] , \mul_b1/fa1_c1[21] ,
         \mul_b1/fa1_c1[20] , \mul_b1/fa1_c1[19] , \mul_b1/fa1_c1[18] ,
         \mul_b1/fa1_c1[17] , \mul_b1/fa1_c1[16] , \mul_b1/fa1_c1[15] ,
         \mul_b1/fa1_c1[14] , \mul_b1/fa1_c1[13] , \mul_b1/fa1_c1[12] ,
         \mul_b1/fa1_c1[11] , \mul_b1/fa1_c1[10] , \mul_b1/fa1_c1[9] ,
         \mul_b1/fa1_c1[8] , \mul_b1/fa1_s1[22] , \mul_b1/fa1_s1[21] ,
         \mul_b1/fa1_s1[20] , \mul_b1/fa1_s1[19] , \mul_b1/fa1_s1[18] ,
         \mul_b1/fa1_s1[17] , \mul_b1/fa1_s1[16] , \mul_b1/fa1_s1[15] ,
         \mul_b1/fa1_s1[14] , \mul_b1/fa1_s1[13] , \mul_b1/fa1_s1[12] ,
         \mul_b1/fa1_s1[11] , \mul_b1/fa1_s1[10] , \mul_b1/fa1_s1[9] ,
         \mul_b1/fa1_s1[8] , \mul_b1/fa1_s1[7] , \mul_b1/fa1_c0[17] ,
         \mul_b1/fa1_c0[16] , \mul_b1/fa1_c0[15] , \mul_b1/fa1_c0[14] ,
         \mul_b1/fa1_c0[13] , \mul_b1/fa1_c0[12] , \mul_b1/fa1_c0[11] ,
         \mul_b1/fa1_c0[10] , \mul_b1/fa1_c0[9] , \mul_b1/fa1_c0[8] ,
         \mul_b1/fa1_c0[7] , \mul_b1/fa1_c0[6] , \mul_b1/fa1_c0[5] ,
         \mul_b1/fa1_c0[4] , \mul_b1/fa1_s0[29] , \mul_b1/fa1_s0[20] ,
         \mul_b1/fa1_s0[19] , \mul_b1/fa1_s0[18] , \mul_b1/fa1_s0[17] ,
         \mul_b1/fa1_s0[16] , \mul_b1/fa1_s0[15] , \mul_b1/fa1_s0[14] ,
         \mul_b1/fa1_s0[13] , \mul_b1/fa1_s0[12] , \mul_b1/fa1_s0[11] ,
         \mul_b1/fa1_s0[10] , \mul_b1/fa1_s0[9] , \mul_b1/fa1_s0[8] ,
         \mul_b1/fa1_s0[7] , \mul_b1/fa1_s0[6] , \mul_b1/fa1_s0[5] ,
         \mul_b1/fa1_s0[4] , \mul_a1/result_sat[15] , \mul_a1/result_sat[14] ,
         \mul_a1/result_sat[13] , \mul_a1/result_sat[12] ,
         \mul_a1/result_sat[11] , \mul_a1/result_sat[10] ,
         \mul_a1/result_sat[9] , \mul_a1/result_sat[8] ,
         \mul_a1/result_sat[7] , \mul_a1/result_sat[6] ,
         \mul_a1/result_sat[5] , \mul_a1/result_sat[4] ,
         \mul_a1/result_sat[3] , \mul_a1/result_sat[2] ,
         \mul_a1/result_sat[1] , \mul_a1/result_sat[0] , \mul_a1/fa1_c2_r[29] ,
         \mul_a1/fa1_c2_r[28] , \mul_a1/fa1_c2_r[27] , \mul_a1/fa1_c2_r[26] ,
         \mul_a1/fa1_c2_r[25] , \mul_a1/fa1_c2_r[24] , \mul_a1/fa1_c2_r[23] ,
         \mul_a1/fa1_c2_r[22] , \mul_a1/fa1_c2_r[21] , \mul_a1/fa1_c2_r[20] ,
         \mul_a1/fa1_c2_r[19] , \mul_a1/fa1_c2_r[18] , \mul_a1/fa1_c2_r[17] ,
         \mul_a1/fa1_c2_r[16] , \mul_a1/fa1_c2_r[15] , \mul_a1/fa1_c2_r[14] ,
         \mul_a1/fa1_s2_r[33] , \mul_a1/fa1_s2_r[32] , \mul_a1/fa1_s2_r[31] ,
         \mul_a1/fa1_s2_r[30] , \mul_a1/fa1_s2_r[29] , \mul_a1/fa1_s2_r[28] ,
         \mul_a1/fa1_s2_r[27] , \mul_a1/fa1_s2_r[26] , \mul_a1/fa1_s2_r[25] ,
         \mul_a1/fa1_s2_r[24] , \mul_a1/fa1_s2_r[23] , \mul_a1/fa1_s2_r[22] ,
         \mul_a1/fa1_s2_r[21] , \mul_a1/fa1_s2_r[20] , \mul_a1/fa1_s2_r[19] ,
         \mul_a1/fa1_s2_r[18] , \mul_a1/fa1_s2_r[17] , \mul_a1/fa1_s2_r[16] ,
         \mul_a1/fa1_s2_r[15] , \mul_a1/fa1_s2_r[14] , \mul_a1/fa1_s2_r[13] ,
         \mul_a1/fa1_c1_r[32] , \mul_a1/fa1_c1_r[31] , \mul_a1/fa1_c1_r[30] ,
         \mul_a1/fa1_c1_r[29] , \mul_a1/fa1_c1_r[28] , \mul_a1/fa1_c1_r[27] ,
         \mul_a1/fa1_c1_r[26] , \mul_a1/fa1_c1_r[25] , \mul_a1/fa1_c1_r[24] ,
         \mul_a1/fa1_c1_r[23] , \mul_a1/fa1_c1_r[22] , \mul_a1/fa1_c1_r[21] ,
         \mul_a1/fa1_c1_r[20] , \mul_a1/fa1_c1_r[19] , \mul_a1/fa1_c1_r[18] ,
         \mul_a1/fa1_c1_r[17] , \mul_a1/fa1_c1_r[16] , \mul_a1/fa1_c1_r[15] ,
         \mul_a1/fa1_c1_r[14] , \mul_a1/fa1_c1_r[13] , \mul_a1/fa1_c1_r[12] ,
         \mul_a1/fa1_c1_r[11] , \mul_a1/fa1_c1_r[10] , \mul_a1/fa1_c1_r[9] ,
         \mul_a1/fa1_c1_r[8] , \mul_a1/fa1_s1_r[33] , \mul_a1/fa1_s1_r[32] ,
         \mul_a1/fa1_s1_r[31] , \mul_a1/fa1_s1_r[30] , \mul_a1/fa1_s1_r[29] ,
         \mul_a1/fa1_s1_r[28] , \mul_a1/fa1_s1_r[27] , \mul_a1/fa1_s1_r[26] ,
         \mul_a1/fa1_s1_r[25] , \mul_a1/fa1_s1_r[24] , \mul_a1/fa1_s1_r[23] ,
         \mul_a1/fa1_s1_r[22] , \mul_a1/fa1_s1_r[21] , \mul_a1/fa1_s1_r[20] ,
         \mul_a1/fa1_s1_r[19] , \mul_a1/fa1_s1_r[18] , \mul_a1/fa1_s1_r[17] ,
         \mul_a1/fa1_s1_r[16] , \mul_a1/fa1_s1_r[15] , \mul_a1/fa1_s1_r[14] ,
         \mul_a1/fa1_s1_r[13] , \mul_a1/fa1_s1_r[12] , \mul_a1/fa1_s1_r[11] ,
         \mul_a1/fa1_s1_r[10] , \mul_a1/fa1_s1_r[9] , \mul_a1/fa1_s1_r[8] ,
         \mul_a1/fa1_s1_r[7] , \mul_a1/fa1_s1_r[6] , \mul_a1/fa1_s0_r[33] ,
         \mul_a1/fa1_s0_r[32] , \mul_a1/fa1_s0_r[31] , \mul_a1/fa1_s0_r[30] ,
         \mul_a1/fa1_s0_r[29] , \mul_a1/fa1_s0_r[28] , \mul_a1/fa1_s0_r[27] ,
         \mul_a1/fa1_s0_r[26] , \mul_a1/fa1_s0_r[25] , \mul_a1/fa1_s0_r[24] ,
         \mul_a1/fa1_s0_r[23] , \mul_a1/fa1_s0_r[22] , \mul_a1/fa1_s0_r[21] ,
         \mul_a1/fa1_s0_r[20] , \mul_a1/fa1_s0_r[19] , \mul_a1/fa1_s0_r[18] ,
         \mul_a1/fa1_s0_r[17] , \mul_a1/fa1_s0_r[16] , \mul_a1/fa1_s0_r[15] ,
         \mul_a1/fa1_s0_r[14] , \mul_a1/fa1_s0_r[13] , \mul_a1/fa1_s0_r[12] ,
         \mul_a1/fa1_s0_r[11] , \mul_a1/fa1_s0_r[10] , \mul_a1/fa1_s0_r[9] ,
         \mul_a1/fa1_s0_r[8] , \mul_a1/fa1_s0_r[7] , \mul_a1/fa1_s0_r[6] ,
         \mul_a1/fa1_c2[29] , \mul_a1/fa1_c2[28] , \mul_a1/fa1_c2[27] ,
         \mul_a1/fa1_c2[26] , \mul_a1/fa1_c2[25] , \mul_a1/fa1_c2[24] ,
         \mul_a1/fa1_c2[23] , \mul_a1/fa1_c2[22] , \mul_a1/fa1_c2[21] ,
         \mul_a1/fa1_c2[20] , \mul_a1/fa1_c2[19] , \mul_a1/fa1_c2[18] ,
         \mul_a1/fa1_c2[17] , \mul_a1/fa1_c2[16] , \mul_a1/fa1_c2[15] ,
         \mul_a1/fa1_c2[14] , \mul_a1/fa1_s2[31] , \mul_a1/fa1_s2[30] ,
         \mul_a1/fa1_s2[29] , \mul_a1/fa1_s2[28] , \mul_a1/fa1_s2[27] ,
         \mul_a1/fa1_s2[26] , \mul_a1/fa1_s2[25] , \mul_a1/fa1_s2[24] ,
         \mul_a1/fa1_s2[23] , \mul_a1/fa1_s2[22] , \mul_a1/fa1_s2[21] ,
         \mul_a1/fa1_s2[20] , \mul_a1/fa1_s2[19] , \mul_a1/fa1_s2[18] ,
         \mul_a1/fa1_s2[17] , \mul_a1/fa1_s2[16] , \mul_a1/fa1_s2[15] ,
         \mul_a1/fa1_s2[14] , \mul_a1/fa1_s2[13] , \mul_a1/fa1_c1[27] ,
         \mul_a1/fa1_c1[22] , \mul_a1/fa1_c1[21] , \mul_a1/fa1_c1[20] ,
         \mul_a1/fa1_c1[19] , \mul_a1/fa1_c1[18] , \mul_a1/fa1_c1[17] ,
         \mul_a1/fa1_c1[16] , \mul_a1/fa1_c1[15] , \mul_a1/fa1_c1[14] ,
         \mul_a1/fa1_c1[13] , \mul_a1/fa1_c1[12] , \mul_a1/fa1_c1[11] ,
         \mul_a1/fa1_c1[10] , \mul_a1/fa1_s1[28] , \mul_a1/fa1_s1[26] ,
         \mul_a1/fa1_s1[25] , \mul_a1/fa1_s1[24] , \mul_a1/fa1_s1[23] ,
         \mul_a1/fa1_s1[22] , \mul_a1/fa1_s1[21] , \mul_a1/fa1_s1[20] ,
         \mul_a1/fa1_s1[19] , \mul_a1/fa1_s1[18] , \mul_a1/fa1_s1[17] ,
         \mul_a1/fa1_s1[16] , \mul_a1/fa1_s1[15] , \mul_a1/fa1_s1[14] ,
         \mul_a1/fa1_s1[13] , \mul_a1/fa1_s1[12] , \mul_a1/fa1_s1[11] ,
         \mul_a1/fa1_s1[10] , \mul_a1/fa1_s1[9] , \mul_a1/fa1_s1[8] ,
         \mul_a1/fa1_s1[7] , n3370, n3371, n3373, n3374, n3376, n3377, n3379,
         n3380, n3382, n3383, n3385, n3386, n3388, n3389, n3391, n3392, n3394,
         n3395, n3397, n3398, n3400, n3401, n3403, n3404, n3406, n3407, n3409,
         n3410, n3412, n3413, n3415, n3416, n3418, n3420, n3422, n3424, n3426,
         n3428, n3430, n3432, n3434, n3436, n3438, n3440, n3442, n3444, n3446,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         \DP_OP_426J1_214_8117/n94 , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056;
  wire   [15:0] x_z1;
  wire   [15:0] x_z2;
  wire   [15:0] y_z1;
  wire   [15:0] p_b0;
  wire   [15:0] p_b1;
  wire   [15:0] p_a1;

  HS65_GS_DFPRQX4 valid_T1_reg ( .D(valid_in), .CP(clk), .RN(rst_n), .Q(
        valid_T1) );
  HS65_GS_DFPRQX4 valid_T2_reg ( .D(valid_T1), .CP(clk), .RN(rst_n), .Q(
        valid_T2) );
  HS65_GS_DFPRQX4 valid_T3_reg ( .D(valid_T2), .CP(clk), .RN(rst_n), .Q(
        valid_T3) );
  HS65_GS_DFPRQX4 valid_out_reg ( .D(valid_T3), .CP(clk), .RN(rst_n), .Q(
        valid_out) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[0]  ( .D(\mul_b0/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[0]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[1]  ( .D(\mul_b0/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[1]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[2]  ( .D(\mul_b0/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[2]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[3]  ( .D(\mul_b0/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[3]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[4]  ( .D(\mul_b0/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[4]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[5]  ( .D(\mul_b0/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[5]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[6]  ( .D(\mul_b0/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[6]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[7]  ( .D(\mul_b0/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[7]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[8]  ( .D(\mul_b0/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[8]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[9]  ( .D(\mul_b0/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[9]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[10]  ( .D(\mul_b0/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[10]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[11]  ( .D(\mul_b0/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[11]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[12]  ( .D(\mul_b0/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[12]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[13]  ( .D(\mul_b0/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[13]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[14]  ( .D(\mul_b0/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[14]) );
  HS65_GS_DFPRQX4 \mul_b0/p_reg[15]  ( .D(\mul_b0/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_b0[15]) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[12]  ( .D(x_z1[0]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[13]  ( .D(x_z1[1]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[14]  ( .D(x_z1[2]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[15]  ( .D(x_z1[3]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[16]  ( .D(x_z1[4]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[17]  ( .D(x_z1[5]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[18]  ( .D(x_z1[6]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[19]  ( .D(x_z1[7]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[20]  ( .D(x_z1[8]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[21]  ( .D(x_z1[9]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[22]  ( .D(x_z1[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[23]  ( .D(x_z1[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[24]  ( .D(x_z1[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[25]  ( .D(x_z1[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[26]  ( .D(x_z1[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[27]  ( .D(n1056), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[28]  ( .D(n1056), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[29]  ( .D(n1056), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[30]  ( .D(n1056), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[31]  ( .D(n1056), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[32]  ( .D(n1056), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s2_r_reg[33]  ( .D(n1056), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[8]  ( .D(x_z1[0]), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[9]  ( .D(x_z1[1]), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[10]  ( .D(x_z1[2]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[11]  ( .D(x_z1[3]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[12]  ( .D(x_z1[4]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[13]  ( .D(x_z1[5]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[14]  ( .D(x_z1[6]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[15]  ( .D(x_z1[7]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[16]  ( .D(x_z1[8]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[17]  ( .D(x_z1[9]), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[18]  ( .D(x_z1[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[19]  ( .D(x_z1[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[20]  ( .D(x_z1[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[21]  ( .D(x_z1[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[22]  ( .D(x_z1[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[23]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[24]  ( .D(n1056), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[25]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[26]  ( .D(n1056), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[27]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[28]  ( .D(n1056), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[29]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[30]  ( .D(n1056), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[31]  ( .D(x_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b0/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[32]  ( .D(n1056), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s1_r_reg[33]  ( .D(n1056), .CP(clk), .RN(rst_n), 
        .Q(\mul_b0/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[5]  ( .D(\mul_b0/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[6]  ( .D(\mul_b0/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[7]  ( .D(\mul_b0/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[8]  ( .D(\mul_b0/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[9]  ( .D(\mul_b0/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[10]  ( .D(\mul_b0/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[11]  ( .D(\mul_b0/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[12]  ( .D(\mul_b0/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[13]  ( .D(\mul_b0/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[14]  ( .D(\mul_b0/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[15]  ( .D(\mul_b0/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[16]  ( .D(\mul_b0/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[17]  ( .D(\mul_b0/fa1_c0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[18]  ( .D(\mul_b0/fa1_c0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[19]  ( .D(\mul_b0/fa1_c0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_c0_r_reg[20]  ( .D(\mul_b0/fa1_c0[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_c0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[6]  ( .D(\mul_b0/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[7]  ( .D(\mul_b0/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[8]  ( .D(\mul_b0/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[9]  ( .D(\mul_b0/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b0/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[10]  ( .D(\mul_b0/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[11]  ( .D(\mul_b0/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[12]  ( .D(\mul_b0/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[13]  ( .D(\mul_b0/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[14]  ( .D(\mul_b0/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[15]  ( .D(\mul_b0/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[16]  ( .D(\mul_b0/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[17]  ( .D(\mul_b0/fa1_s0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[18]  ( .D(\mul_b0/fa1_s0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[19]  ( .D(\mul_b0/fa1_s0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[20]  ( .D(\mul_b0/fa1_s0[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[21]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[22]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[23]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[24]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[25]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[26]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[27]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[28]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[29]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[30]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[31]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[32]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b0/fa1_s0_r_reg[33]  ( .D(\mul_b0/fa1_s0[30] ), .CP(clk), .RN(rst_n), .Q(\mul_b0/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[0]  ( .D(\mul_b1/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[0]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[1]  ( .D(\mul_b1/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[1]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[2]  ( .D(\mul_b1/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[2]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[3]  ( .D(\mul_b1/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[3]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[4]  ( .D(\mul_b1/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[4]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[5]  ( .D(\mul_b1/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[5]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[6]  ( .D(\mul_b1/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[6]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[7]  ( .D(\mul_b1/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[7]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[8]  ( .D(\mul_b1/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[8]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[9]  ( .D(\mul_b1/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[9]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[10]  ( .D(\mul_b1/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[10]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[11]  ( .D(\mul_b1/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[11]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[12]  ( .D(\mul_b1/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[12]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[13]  ( .D(\mul_b1/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[13]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[14]  ( .D(\mul_b1/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[14]) );
  HS65_GS_DFPRQX4 \mul_b1/p_reg[15]  ( .D(\mul_b1/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_b1[15]) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[12]  ( .D(\mul_b1/fa1_s1[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s2_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[13]  ( .D(x_z2[1]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[14]  ( .D(x_z2[2]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[15]  ( .D(x_z2[3]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[16]  ( .D(x_z2[4]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[17]  ( .D(x_z2[5]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[18]  ( .D(x_z2[6]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[19]  ( .D(x_z2[7]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[20]  ( .D(x_z2[8]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[21]  ( .D(x_z2[9]), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[22]  ( .D(x_z2[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[23]  ( .D(x_z2[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[24]  ( .D(x_z2[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[25]  ( .D(x_z2[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[26]  ( .D(x_z2[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[27]  ( .D(n1055), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[28]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[29]  ( .D(n1055), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[30]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[31]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[32]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s2_r_reg[33]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[8]  ( .D(\mul_b1/fa1_c1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[9]  ( .D(\mul_b1/fa1_c1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[10]  ( .D(\mul_b1/fa1_c1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[11]  ( .D(\mul_b1/fa1_c1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[12]  ( .D(\mul_b1/fa1_c1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[13]  ( .D(\mul_b1/fa1_c1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[14]  ( .D(\mul_b1/fa1_c1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[15]  ( .D(\mul_b1/fa1_c1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[16]  ( .D(\mul_b1/fa1_c1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[17]  ( .D(\mul_b1/fa1_c1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[18]  ( .D(\mul_b1/fa1_c1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[19]  ( .D(\mul_b1/fa1_c1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[20]  ( .D(\mul_b1/fa1_c1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[21]  ( .D(\mul_b1/fa1_c1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[22]  ( .D(\mul_b1/fa1_c1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[23]  ( .D(x_z2[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_b1/fa1_c1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[24]  ( .D(n1055), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[25]  ( .D(n1055), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[26]  ( .D(n1055), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[27]  ( .D(n1055), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[28]  ( .D(n1055), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[29]  ( .D(n1055), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[30]  ( .D(n1055), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[31]  ( .D(n1055), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c1_r_reg[32]  ( .D(n1055), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[7]  ( .D(\mul_b1/fa1_s1[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s1_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[8]  ( .D(\mul_b1/fa1_s1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[9]  ( .D(\mul_b1/fa1_s1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[10]  ( .D(\mul_b1/fa1_s1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[11]  ( .D(\mul_b1/fa1_s1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[12]  ( .D(\mul_b1/fa1_s1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[13]  ( .D(\mul_b1/fa1_s1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[14]  ( .D(\mul_b1/fa1_s1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[15]  ( .D(\mul_b1/fa1_s1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[16]  ( .D(\mul_b1/fa1_s1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[17]  ( .D(\mul_b1/fa1_s1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[18]  ( .D(\mul_b1/fa1_s1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[19]  ( .D(\mul_b1/fa1_s1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[20]  ( .D(\mul_b1/fa1_s1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[21]  ( .D(\mul_b1/fa1_s1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s1_r_reg[22]  ( .D(\mul_b1/fa1_s1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[3]  ( .D(n1053), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[3] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[4]  ( .D(\mul_b1/fa1_c0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[5]  ( .D(\mul_b1/fa1_c0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[6]  ( .D(\mul_b1/fa1_c0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[7]  ( .D(\mul_b1/fa1_c0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[8]  ( .D(\mul_b1/fa1_c0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[9]  ( .D(\mul_b1/fa1_c0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_c0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[10]  ( .D(\mul_b1/fa1_c0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[11]  ( .D(\mul_b1/fa1_c0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[12]  ( .D(\mul_b1/fa1_c0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[13]  ( .D(\mul_b1/fa1_c0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[14]  ( .D(\mul_b1/fa1_c0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[15]  ( .D(\mul_b1/fa1_c0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[16]  ( .D(\mul_b1/fa1_c0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[17]  ( .D(\mul_b1/fa1_c0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_c0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[18]  ( .D(n578), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[19]  ( .D(n580), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[20]  ( .D(n1051), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[21]  ( .D(n1051), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[22]  ( .D(n1051), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[23]  ( .D(n1051), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[24]  ( .D(n1051), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[25]  ( .D(n1051), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[26]  ( .D(n1051), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[27]  ( .D(n1051), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[28]  ( .D(n1051), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[29]  ( .D(n1051), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[30]  ( .D(n1051), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[31]  ( .D(n1051), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_c0_r_reg[32]  ( .D(n1051), .CP(clk), .RN(rst_n), 
        .Q(\mul_b1/fa1_c0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[4]  ( .D(\mul_b1/fa1_s0[4] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[4] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[5]  ( .D(\mul_b1/fa1_s0[5] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[5] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[6]  ( .D(\mul_b1/fa1_s0[6] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[7]  ( .D(\mul_b1/fa1_s0[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[8]  ( .D(\mul_b1/fa1_s0[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[9]  ( .D(\mul_b1/fa1_s0[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_b1/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[10]  ( .D(\mul_b1/fa1_s0[10] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[11]  ( .D(\mul_b1/fa1_s0[11] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[12]  ( .D(\mul_b1/fa1_s0[12] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[13]  ( .D(\mul_b1/fa1_s0[13] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[14]  ( .D(\mul_b1/fa1_s0[14] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[15]  ( .D(\mul_b1/fa1_s0[15] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[16]  ( .D(\mul_b1/fa1_s0[16] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[17]  ( .D(\mul_b1/fa1_s0[17] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[18]  ( .D(\mul_b1/fa1_s0[18] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[19]  ( .D(\mul_b1/fa1_s0[19] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[20]  ( .D(\mul_b1/fa1_s0[20] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[21]  ( .D(\mul_b1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[22]  ( .D(\mul_b1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[23]  ( .D(\mul_b1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[24]  ( .D(\mul_b1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[25]  ( .D(\mul_b1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[26]  ( .D(\mul_b1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[27]  ( .D(\mul_b1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[28]  ( .D(\mul_b1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[29]  ( .D(\mul_b1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[30]  ( .D(\mul_b1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[31]  ( .D(\mul_b1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[32]  ( .D(\mul_b1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_b1/fa1_s0_r_reg[33]  ( .D(\mul_b1/fa1_s0[29] ), .CP(clk), .RN(rst_n), .Q(\mul_b1/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[0]  ( .D(\mul_a1/result_sat[0] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[0]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[1]  ( .D(\mul_a1/result_sat[1] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[1]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[2]  ( .D(\mul_a1/result_sat[2] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[2]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[3]  ( .D(\mul_a1/result_sat[3] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[3]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[4]  ( .D(\mul_a1/result_sat[4] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[4]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[5]  ( .D(\mul_a1/result_sat[5] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[5]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[6]  ( .D(\mul_a1/result_sat[6] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[6]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[7]  ( .D(\mul_a1/result_sat[7] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[7]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[8]  ( .D(\mul_a1/result_sat[8] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[8]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[9]  ( .D(\mul_a1/result_sat[9] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[9]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[10]  ( .D(\mul_a1/result_sat[10] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[10]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[11]  ( .D(\mul_a1/result_sat[11] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[11]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[12]  ( .D(\mul_a1/result_sat[12] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[12]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[13]  ( .D(\mul_a1/result_sat[13] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[13]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[14]  ( .D(\mul_a1/result_sat[14] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[14]) );
  HS65_GS_DFPRQX4 \mul_a1/p_reg[15]  ( .D(\mul_a1/result_sat[15] ), .CP(clk), 
        .RN(rst_n), .Q(p_a1[15]) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[13]  ( .D(\mul_a1/fa1_s2[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[14]  ( .D(\mul_a1/fa1_s2[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[15]  ( .D(\mul_a1/fa1_s2[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[16]  ( .D(\mul_a1/fa1_s2[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[17]  ( .D(\mul_a1/fa1_s2[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[18]  ( .D(\mul_a1/fa1_s2[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[19]  ( .D(\mul_a1/fa1_s2[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[20]  ( .D(\mul_a1/fa1_s2[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[21]  ( .D(\mul_a1/fa1_s2[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[22]  ( .D(\mul_a1/fa1_s2[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[23]  ( .D(\mul_a1/fa1_s2[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[24]  ( .D(\mul_a1/fa1_s2[24] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[25]  ( .D(\mul_a1/fa1_s2[25] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[26]  ( .D(\mul_a1/fa1_s2[26] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[27]  ( .D(\mul_a1/fa1_s2[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[28]  ( .D(\mul_a1/fa1_s2[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[29]  ( .D(\mul_a1/fa1_s2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[30]  ( .D(\mul_a1/fa1_s2[30] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[31]  ( .D(\mul_a1/fa1_s2[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[32]  ( .D(\mul_a1/fa1_s2[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s2_r_reg[33]  ( .D(\mul_a1/fa1_s2[31] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s2_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[8]  ( .D(n1049), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_c1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[9]  ( .D(n1050), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_c1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[10]  ( .D(\mul_a1/fa1_c1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[11]  ( .D(\mul_a1/fa1_c1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[12]  ( .D(\mul_a1/fa1_c1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[13]  ( .D(\mul_a1/fa1_c1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[14]  ( .D(\mul_a1/fa1_c1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[15]  ( .D(\mul_a1/fa1_c1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[16]  ( .D(\mul_a1/fa1_c1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[17]  ( .D(\mul_a1/fa1_c1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[18]  ( .D(\mul_a1/fa1_c1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[19]  ( .D(\mul_a1/fa1_c1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[20]  ( .D(\mul_a1/fa1_c1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[21]  ( .D(\mul_a1/fa1_c1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[22]  ( .D(\mul_a1/fa1_c1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[23]  ( .D(n463), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_c1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[24]  ( .D(n465), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_c1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[25]  ( .D(n1054), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_c1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[26]  ( .D(n1052), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_c1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[27]  ( .D(\mul_a1/fa1_c1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[28]  ( .D(\mul_a1/fa1_c1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[29]  ( .D(\mul_a1/fa1_c1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[30]  ( .D(\mul_a1/fa1_c1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[31]  ( .D(\mul_a1/fa1_c1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c1_r_reg[32]  ( .D(\mul_a1/fa1_c1[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[6]  ( .D(\mul_a1/fa1_s2[13] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[6] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[7]  ( .D(\mul_a1/fa1_s1[7] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[8]  ( .D(\mul_a1/fa1_s1[8] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[9]  ( .D(\mul_a1/fa1_s1[9] ), .CP(clk), 
        .RN(rst_n), .Q(\mul_a1/fa1_s1_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[10]  ( .D(\mul_a1/fa1_s1[10] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[11]  ( .D(\mul_a1/fa1_s1[11] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[12]  ( .D(\mul_a1/fa1_s1[12] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[13]  ( .D(\mul_a1/fa1_s1[13] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[14]  ( .D(\mul_a1/fa1_s1[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[15]  ( .D(\mul_a1/fa1_s1[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[16]  ( .D(\mul_a1/fa1_s1[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[17]  ( .D(\mul_a1/fa1_s1[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[18]  ( .D(\mul_a1/fa1_s1[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[19]  ( .D(\mul_a1/fa1_s1[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[20]  ( .D(\mul_a1/fa1_s1[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[21]  ( .D(\mul_a1/fa1_s1[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[22]  ( .D(\mul_a1/fa1_s1[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[23]  ( .D(\mul_a1/fa1_s1[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[24]  ( .D(\mul_a1/fa1_s1[24] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[25]  ( .D(\mul_a1/fa1_s1[25] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[26]  ( .D(\mul_a1/fa1_s1[26] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[27]  ( .D(\mul_a1/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[28]  ( .D(\mul_a1/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[29]  ( .D(\mul_a1/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[30]  ( .D(\mul_a1/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[31]  ( .D(\mul_a1/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[32]  ( .D(\mul_a1/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s1_r_reg[33]  ( .D(\mul_a1/fa1_s1[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s1_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[6]  ( .D(y_z1[2]), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[6] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[7]  ( .D(y_z1[3]), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[7] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[8]  ( .D(y_z1[4]), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[8] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[9]  ( .D(y_z1[5]), .CP(clk), .RN(rst_n), 
        .Q(\mul_a1/fa1_s0_r[9] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[10]  ( .D(y_z1[6]), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[10] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[11]  ( .D(y_z1[7]), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[11] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[12]  ( .D(y_z1[8]), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[12] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[13]  ( .D(y_z1[9]), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[13] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[14]  ( .D(y_z1[10]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[15]  ( .D(y_z1[11]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[16]  ( .D(y_z1[12]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[17]  ( .D(y_z1[13]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[18]  ( .D(y_z1[14]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[19]  ( .D(\DP_OP_426J1_214_8117/n94 ), 
        .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[20]  ( .D(\DP_OP_426J1_214_8117/n94 ), 
        .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[21]  ( .D(\DP_OP_426J1_214_8117/n94 ), 
        .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[22]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[23]  ( .D(\DP_OP_426J1_214_8117/n94 ), 
        .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_s0_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[24]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[25]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[26]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[27]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[28]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[29]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[29] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[30]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[30] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[31]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[31] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[32]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[32] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_s0_r_reg[33]  ( .D(y_z1[15]), .CP(clk), .RN(
        rst_n), .Q(\mul_a1/fa1_s0_r[33] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[14]  ( .D(\mul_a1/fa1_c2[14] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[14] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[15]  ( .D(\mul_a1/fa1_c2[15] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[15] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[16]  ( .D(\mul_a1/fa1_c2[16] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[16] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[17]  ( .D(\mul_a1/fa1_c2[17] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[17] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[18]  ( .D(\mul_a1/fa1_c2[18] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[18] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[19]  ( .D(\mul_a1/fa1_c2[19] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[19] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[20]  ( .D(\mul_a1/fa1_c2[20] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[20] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[21]  ( .D(\mul_a1/fa1_c2[21] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[21] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[22]  ( .D(\mul_a1/fa1_c2[22] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[22] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[23]  ( .D(\mul_a1/fa1_c2[23] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[23] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[24]  ( .D(\mul_a1/fa1_c2[24] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[24] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[25]  ( .D(\mul_a1/fa1_c2[25] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[25] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[26]  ( .D(\mul_a1/fa1_c2[26] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[26] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[27]  ( .D(\mul_a1/fa1_c2[27] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[27] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[28]  ( .D(\mul_a1/fa1_c2[28] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[28] ) );
  HS65_GS_DFPRQX4 \mul_a1/fa1_c2_r_reg[29]  ( .D(\mul_a1/fa1_c2[29] ), .CP(clk), .RN(rst_n), .Q(\mul_a1/fa1_c2_r[29] ) );
  HS65_GS_DFPRQX4 \x_z1_reg[15]  ( .D(n3464), .CP(clk), .RN(rst_n), .Q(
        x_z1[15]) );
  HS65_GS_DFPRQX4 \x_z1_reg[14]  ( .D(n3463), .CP(clk), .RN(rst_n), .Q(
        x_z1[14]) );
  HS65_GS_DFPRQX4 \x_z1_reg[13]  ( .D(n3462), .CP(clk), .RN(rst_n), .Q(
        x_z1[13]) );
  HS65_GS_DFPRQX4 \x_z1_reg[12]  ( .D(n3461), .CP(clk), .RN(rst_n), .Q(
        x_z1[12]) );
  HS65_GS_DFPRQX4 \x_z1_reg[11]  ( .D(n3460), .CP(clk), .RN(rst_n), .Q(
        x_z1[11]) );
  HS65_GS_DFPRQX4 \x_z1_reg[10]  ( .D(n3459), .CP(clk), .RN(rst_n), .Q(
        x_z1[10]) );
  HS65_GS_DFPRQX4 \x_z1_reg[9]  ( .D(n3458), .CP(clk), .RN(rst_n), .Q(x_z1[9])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[8]  ( .D(n3457), .CP(clk), .RN(rst_n), .Q(x_z1[8])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[7]  ( .D(n3456), .CP(clk), .RN(rst_n), .Q(x_z1[7])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[6]  ( .D(n3455), .CP(clk), .RN(rst_n), .Q(x_z1[6])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[5]  ( .D(n3454), .CP(clk), .RN(rst_n), .Q(x_z1[5])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[4]  ( .D(n3453), .CP(clk), .RN(rst_n), .Q(x_z1[4])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[3]  ( .D(n3452), .CP(clk), .RN(rst_n), .Q(x_z1[3])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[2]  ( .D(n3451), .CP(clk), .RN(rst_n), .Q(x_z1[2])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[1]  ( .D(n3450), .CP(clk), .RN(rst_n), .Q(x_z1[1])
         );
  HS65_GS_DFPRQX4 \x_z1_reg[0]  ( .D(n3449), .CP(clk), .RN(rst_n), .Q(x_z1[0])
         );
  HS65_GS_DFPRQX4 \x_z2_reg[15]  ( .D(n3448), .CP(clk), .RN(rst_n), .Q(
        x_z2[15]) );
  HS65_GS_DFPRQX4 \x_z2_reg[14]  ( .D(n3446), .CP(clk), .RN(rst_n), .Q(
        x_z2[14]) );
  HS65_GS_DFPRQX4 \x_z2_reg[13]  ( .D(n3444), .CP(clk), .RN(rst_n), .Q(
        x_z2[13]) );
  HS65_GS_DFPRQX4 \x_z2_reg[12]  ( .D(n3442), .CP(clk), .RN(rst_n), .Q(
        x_z2[12]) );
  HS65_GS_DFPRQX4 \x_z2_reg[11]  ( .D(n3440), .CP(clk), .RN(rst_n), .Q(
        x_z2[11]) );
  HS65_GS_DFPRQX4 \x_z2_reg[10]  ( .D(n3438), .CP(clk), .RN(rst_n), .Q(
        x_z2[10]) );
  HS65_GS_DFPRQX4 \x_z2_reg[9]  ( .D(n3436), .CP(clk), .RN(rst_n), .Q(x_z2[9])
         );
  HS65_GS_DFPRQX4 \x_z2_reg[8]  ( .D(n3434), .CP(clk), .RN(rst_n), .Q(x_z2[8])
         );
  HS65_GS_DFPRQX4 \x_z2_reg[7]  ( .D(n3432), .CP(clk), .RN(rst_n), .Q(x_z2[7])
         );
  HS65_GS_DFPRQX4 \x_z2_reg[6]  ( .D(n3430), .CP(clk), .RN(rst_n), .Q(x_z2[6])
         );
  HS65_GS_DFPRQX4 \x_z2_reg[5]  ( .D(n3428), .CP(clk), .RN(rst_n), .Q(x_z2[5])
         );
  HS65_GS_DFPRQX4 \x_z2_reg[4]  ( .D(n3426), .CP(clk), .RN(rst_n), .Q(x_z2[4])
         );
  HS65_GS_DFPRQX4 \x_z2_reg[3]  ( .D(n3424), .CP(clk), .RN(rst_n), .Q(x_z2[3])
         );
  HS65_GS_DFPRQX4 \x_z2_reg[2]  ( .D(n3422), .CP(clk), .RN(rst_n), .Q(x_z2[2])
         );
  HS65_GS_DFPRQX4 \x_z2_reg[1]  ( .D(n3420), .CP(clk), .RN(rst_n), .Q(x_z2[1])
         );
  HS65_GS_DFPRQX4 \x_z2_reg[0]  ( .D(n3418), .CP(clk), .RN(rst_n), .Q(
        \mul_b1/fa1_s1[7] ) );
  HS65_GS_DFPRQX4 \data_out_reg[15]  ( .D(n3416), .CP(clk), .RN(rst_n), .Q(
        data_out[15]) );
  HS65_GS_DFPRQX4 \y_z1_reg[15]  ( .D(n3415), .CP(clk), .RN(rst_n), .Q(
        y_z1[15]) );
  HS65_GS_DFPRQX4 \data_out_reg[14]  ( .D(n3413), .CP(clk), .RN(rst_n), .Q(
        data_out[14]) );
  HS65_GS_DFPRQX4 \y_z1_reg[14]  ( .D(n3412), .CP(clk), .RN(rst_n), .Q(
        y_z1[14]) );
  HS65_GS_DFPRQX4 \data_out_reg[13]  ( .D(n3410), .CP(clk), .RN(rst_n), .Q(
        data_out[13]) );
  HS65_GS_DFPRQX4 \y_z1_reg[13]  ( .D(n3409), .CP(clk), .RN(rst_n), .Q(
        y_z1[13]) );
  HS65_GS_DFPRQX4 \data_out_reg[12]  ( .D(n3407), .CP(clk), .RN(rst_n), .Q(
        data_out[12]) );
  HS65_GS_DFPRQX4 \y_z1_reg[12]  ( .D(n3406), .CP(clk), .RN(rst_n), .Q(
        y_z1[12]) );
  HS65_GS_DFPRQX4 \data_out_reg[11]  ( .D(n3404), .CP(clk), .RN(rst_n), .Q(
        data_out[11]) );
  HS65_GS_DFPRQX4 \y_z1_reg[11]  ( .D(n3403), .CP(clk), .RN(rst_n), .Q(
        y_z1[11]) );
  HS65_GS_DFPRQX4 \data_out_reg[10]  ( .D(n3401), .CP(clk), .RN(rst_n), .Q(
        data_out[10]) );
  HS65_GS_DFPRQX4 \y_z1_reg[10]  ( .D(n3400), .CP(clk), .RN(rst_n), .Q(
        y_z1[10]) );
  HS65_GS_DFPRQX4 \data_out_reg[9]  ( .D(n3398), .CP(clk), .RN(rst_n), .Q(
        data_out[9]) );
  HS65_GS_DFPRQX4 \y_z1_reg[9]  ( .D(n3397), .CP(clk), .RN(rst_n), .Q(y_z1[9])
         );
  HS65_GS_DFPRQX4 \data_out_reg[8]  ( .D(n3395), .CP(clk), .RN(rst_n), .Q(
        data_out[8]) );
  HS65_GS_DFPRQX4 \y_z1_reg[8]  ( .D(n3394), .CP(clk), .RN(rst_n), .Q(y_z1[8])
         );
  HS65_GS_DFPRQX4 \data_out_reg[7]  ( .D(n3392), .CP(clk), .RN(rst_n), .Q(
        data_out[7]) );
  HS65_GS_DFPRQX4 \y_z1_reg[7]  ( .D(n3391), .CP(clk), .RN(rst_n), .Q(y_z1[7])
         );
  HS65_GS_DFPRQX4 \data_out_reg[6]  ( .D(n3389), .CP(clk), .RN(rst_n), .Q(
        data_out[6]) );
  HS65_GS_DFPRQX4 \y_z1_reg[6]  ( .D(n3388), .CP(clk), .RN(rst_n), .Q(y_z1[6])
         );
  HS65_GS_DFPRQX4 \data_out_reg[5]  ( .D(n3386), .CP(clk), .RN(rst_n), .Q(
        data_out[5]) );
  HS65_GS_DFPRQX4 \y_z1_reg[5]  ( .D(n3385), .CP(clk), .RN(rst_n), .Q(y_z1[5])
         );
  HS65_GS_DFPRQX4 \data_out_reg[4]  ( .D(n3383), .CP(clk), .RN(rst_n), .Q(
        data_out[4]) );
  HS65_GS_DFPRQX4 \y_z1_reg[4]  ( .D(n3382), .CP(clk), .RN(rst_n), .Q(y_z1[4])
         );
  HS65_GS_DFPRQX4 \data_out_reg[3]  ( .D(n3380), .CP(clk), .RN(rst_n), .Q(
        data_out[3]) );
  HS65_GS_DFPRQX4 \y_z1_reg[3]  ( .D(n3379), .CP(clk), .RN(rst_n), .Q(y_z1[3])
         );
  HS65_GS_DFPRQX4 \data_out_reg[2]  ( .D(n3377), .CP(clk), .RN(rst_n), .Q(
        data_out[2]) );
  HS65_GS_DFPRQX4 \y_z1_reg[2]  ( .D(n3376), .CP(clk), .RN(rst_n), .Q(y_z1[2])
         );
  HS65_GS_DFPRQX4 \data_out_reg[1]  ( .D(n3374), .CP(clk), .RN(rst_n), .Q(
        data_out[1]) );
  HS65_GS_DFPRQX4 \y_z1_reg[1]  ( .D(n3373), .CP(clk), .RN(rst_n), .Q(y_z1[1])
         );
  HS65_GS_DFPRQX4 \data_out_reg[0]  ( .D(n3371), .CP(clk), .RN(rst_n), .Q(
        data_out[0]) );
  HS65_GS_DFPRQX4 \y_z1_reg[0]  ( .D(n3370), .CP(clk), .RN(rst_n), .Q(
        \mul_a1/fa1_s2[13] ) );
  HS65_GS_AND2X4 U3 ( .A(\mul_b0/fa1_s0_r[28] ), .B(\mul_b0/fa1_s1_r[28] ), 
        .Z(n2) );
  HS65_GSS_XOR2X3 U4 ( .A(\mul_b0/fa1_s0_r[29] ), .B(\mul_b0/fa1_s1_r[29] ), 
        .Z(n1) );
  HS65_GS_AND2X4 U5 ( .A(\mul_b0/fa1_s1_r[29] ), .B(\mul_b0/fa1_s0_r[29] ), 
        .Z(n69) );
  HS65_GSS_XOR2X3 U6 ( .A(\mul_b0/fa1_s0_r[30] ), .B(\mul_b0/fa1_s1_r[30] ), 
        .Z(n68) );
  HS65_GS_AND2X4 U7 ( .A(\mul_b0/fa1_s1_r[27] ), .B(\mul_b0/fa1_s0_r[27] ), 
        .Z(n66) );
  HS65_GSS_XOR2X3 U8 ( .A(\mul_b0/fa1_s0_r[28] ), .B(\mul_b0/fa1_s1_r[28] ), 
        .Z(n65) );
  HS65_GS_FA1X4 U9 ( .A0(\mul_b0/fa1_s2_r[29] ), .B0(n2), .CI(n1), .CO(n531), 
        .S0(n533) );
  HS65_GS_AND2X4 U10 ( .A(\mul_b0/fa1_s0_r[23] ), .B(\mul_b0/fa1_s1_r[23] ), 
        .Z(n4) );
  HS65_GSS_XOR2X3 U11 ( .A(\mul_b0/fa1_s0_r[24] ), .B(\mul_b0/fa1_s1_r[24] ), 
        .Z(n3) );
  HS65_GS_AND2X4 U12 ( .A(\mul_b0/fa1_s1_r[24] ), .B(\mul_b0/fa1_s0_r[24] ), 
        .Z(n60) );
  HS65_GSS_XOR2X3 U13 ( .A(\mul_b0/fa1_s0_r[25] ), .B(\mul_b0/fa1_s1_r[25] ), 
        .Z(n59) );
  HS65_GS_FA1X4 U14 ( .A0(\mul_b0/fa1_s2_r[24] ), .B0(n4), .CI(n3), .CO(n819), 
        .S0(n815) );
  HS65_GSS_XOR2X3 U15 ( .A(\mul_b0/fa1_s0_r[23] ), .B(\mul_b0/fa1_s1_r[23] ), 
        .Z(n58) );
  HS65_GS_AND2X4 U16 ( .A(\mul_b0/fa1_s1_r[22] ), .B(\mul_b0/fa1_s0_r[22] ), 
        .Z(n57) );
  HS65_GS_FA1X4 U17 ( .A0(\mul_b0/fa1_s0_r[20] ), .B0(\mul_b0/fa1_s1_r[20] ), 
        .CI(\mul_b0/fa1_c0_r[19] ), .CO(n54), .S0(n5) );
  HS65_GS_FA1X4 U18 ( .A0(\mul_b0/fa1_s0_r[19] ), .B0(\mul_b0/fa1_s1_r[19] ), 
        .CI(\mul_b0/fa1_c0_r[18] ), .CO(n6), .S0(n7) );
  HS65_GS_FA1X4 U19 ( .A0(\mul_b0/fa1_s2_r[20] ), .B0(n6), .CI(n5), .CO(n803), 
        .S0(n798) );
  HS65_GS_FA1X4 U20 ( .A0(\mul_b0/fa1_s0_r[18] ), .B0(\mul_b0/fa1_s1_r[18] ), 
        .CI(\mul_b0/fa1_c0_r[17] ), .CO(n8), .S0(n51) );
  HS65_GS_FA1X4 U21 ( .A0(\mul_b0/fa1_s2_r[19] ), .B0(n8), .CI(n7), .CO(n799), 
        .S0(n794) );
  HS65_GS_FA1X4 U22 ( .A0(\mul_b0/fa1_s0_r[15] ), .B0(\mul_b0/fa1_s1_r[15] ), 
        .CI(\mul_b0/fa1_c0_r[14] ), .CO(n45), .S0(n10) );
  HS65_GS_FA1X4 U23 ( .A0(\mul_b0/fa1_s0_r[14] ), .B0(\mul_b0/fa1_s1_r[14] ), 
        .CI(\mul_b0/fa1_c0_r[13] ), .CO(n9), .S0(n12) );
  HS65_GS_FA1X4 U24 ( .A0(\mul_b0/fa1_s0_r[13] ), .B0(\mul_b0/fa1_s1_r[13] ), 
        .CI(\mul_b0/fa1_c0_r[12] ), .CO(n11), .S0(n13) );
  HS65_GS_FA1X4 U25 ( .A0(\mul_b0/fa1_s2_r[15] ), .B0(n10), .CI(n9), .CO(n572), 
        .S0(n42) );
  HS65_GS_FA1X4 U26 ( .A0(\mul_b0/fa1_s2_r[14] ), .B0(n12), .CI(n11), .CO(n41), 
        .S0(n38) );
  HS65_GSS_XNOR2X3 U27 ( .A(n42), .B(n41), .Z(n1041) );
  HS65_GS_IVX2 U28 ( .A(n1041), .Z(n40) );
  HS65_GS_AOI12X2 U29 ( .A(n37), .B(n38), .C(n40), .Z(n1040) );
  HS65_GS_NAND2X2 U30 ( .A(n38), .B(n37), .Z(n36) );
  HS65_GS_IVX2 U31 ( .A(n36), .Z(n39) );
  HS65_GS_FA1X4 U32 ( .A0(\mul_b0/fa1_s2_r[13] ), .B0(n14), .CI(n13), .CO(n37), 
        .S0(n35) );
  HS65_GS_FA1X4 U33 ( .A0(\mul_b0/fa1_s0_r[12] ), .B0(\mul_b0/fa1_s1_r[12] ), 
        .CI(\mul_b0/fa1_c0_r[11] ), .CO(n14), .S0(n15) );
  HS65_GS_FA1X4 U34 ( .A0(\mul_b0/fa1_s2_r[12] ), .B0(n16), .CI(n15), .CO(n34), 
        .S0(n32) );
  HS65_GS_FA1X4 U35 ( .A0(\mul_b0/fa1_s0_r[11] ), .B0(\mul_b0/fa1_s1_r[11] ), 
        .CI(\mul_b0/fa1_c0_r[10] ), .CO(n16), .S0(n29) );
  HS65_GS_FA1X4 U36 ( .A0(\mul_b0/fa1_s0_r[10] ), .B0(\mul_b0/fa1_s1_r[10] ), 
        .CI(\mul_b0/fa1_c0_r[9] ), .CO(n30), .S0(n26) );
  HS65_GS_NOR2X2 U37 ( .A(n27), .B(n26), .Z(n24) );
  HS65_GS_FA1X4 U38 ( .A0(\mul_b0/fa1_s0_r[8] ), .B0(\mul_b0/fa1_s1_r[8] ), 
        .CI(\mul_b0/fa1_c0_r[7] ), .CO(n22), .S0(n19) );
  HS65_GS_AND2X4 U39 ( .A(\mul_b0/fa1_c0_r[5] ), .B(\mul_b0/fa1_s0_r[6] ), .Z(
        n17) );
  HS65_GS_PAOI2X1 U40 ( .A(\mul_b0/fa1_s0_r[7] ), .B(\mul_b0/fa1_c0_r[6] ), 
        .P(n17), .Z(n18) );
  HS65_GS_NOR2AX3 U41 ( .A(n19), .B(n18), .Z(n21) );
  HS65_GS_FA1X4 U42 ( .A0(\mul_b0/fa1_s0_r[9] ), .B0(\mul_b0/fa1_s1_r[9] ), 
        .CI(\mul_b0/fa1_c0_r[8] ), .CO(n27), .S0(n20) );
  HS65_GS_PAOI2X1 U43 ( .A(n22), .B(n21), .P(n20), .Z(n23) );
  HS65_GS_NOR2X2 U44 ( .A(n24), .B(n23), .Z(n25) );
  HS65_GS_AO12X4 U45 ( .A(n27), .B(n26), .C(n25), .Z(n28) );
  HS65_GS_PAOI2X1 U46 ( .A(n30), .B(n29), .P(n28), .Z(n31) );
  HS65_GS_NOR2AX3 U47 ( .A(n32), .B(n31), .Z(n33) );
  HS65_GS_PAOI2X1 U48 ( .A(n35), .B(n34), .P(n33), .Z(n595) );
  HS65_GS_OAI21X2 U49 ( .A(n38), .B(n37), .C(n36), .Z(n594) );
  HS65_GS_NOR2X2 U50 ( .A(n595), .B(n594), .Z(n1042) );
  HS65_GS_AOI12X2 U51 ( .A(n40), .B(n39), .C(n1042), .Z(n1044) );
  HS65_GS_NAND2X2 U52 ( .A(n42), .B(n41), .Z(n43) );
  HS65_GS_OAI21X2 U53 ( .A(n1040), .B(n1044), .C(n43), .Z(n574) );
  HS65_GS_PAOI2X1 U54 ( .A(n572), .B(n573), .P(n574), .Z(n546) );
  HS65_GS_FA1X4 U55 ( .A0(\mul_b0/fa1_s0_r[16] ), .B0(\mul_b0/fa1_s1_r[16] ), 
        .CI(\mul_b0/fa1_c0_r[15] ), .CO(n50), .S0(n44) );
  HS65_GS_FA1X4 U56 ( .A0(\mul_b0/fa1_s0_r[17] ), .B0(\mul_b0/fa1_s1_r[17] ), 
        .CI(\mul_b0/fa1_c0_r[16] ), .CO(n52), .S0(n49) );
  HS65_GS_FA1X4 U57 ( .A0(\mul_b0/fa1_s2_r[16] ), .B0(n45), .CI(n44), .CO(n46), 
        .S0(n573) );
  HS65_GS_NAND2X2 U58 ( .A(n47), .B(n46), .Z(n48) );
  HS65_GS_OAI21X2 U59 ( .A(n47), .B(n46), .C(n48), .Z(n545) );
  HS65_GS_OAI21X2 U60 ( .A(n546), .B(n545), .C(n48), .Z(n791) );
  HS65_GS_FA1X4 U61 ( .A0(\mul_b0/fa1_s2_r[17] ), .B0(n50), .CI(n49), .CO(n790), .S0(n47) );
  HS65_GS_FA1X4 U62 ( .A0(\mul_b0/fa1_s2_r[18] ), .B0(n52), .CI(n51), .CO(n795), .S0(n789) );
  HS65_GS_FA1X4 U63 ( .A0(\mul_b0/fa1_s2_r[21] ), .B0(n54), .CI(n53), .CO(n806), .S0(n802) );
  HS65_GS_FA1X4 U64 ( .A0(\mul_b0/fa1_s0_r[21] ), .B0(\mul_b0/fa1_s1_r[21] ), 
        .CI(\mul_b0/fa1_c0_r[20] ), .CO(n56), .S0(n53) );
  HS65_GSS_XOR2X3 U65 ( .A(\mul_b0/fa1_s0_r[22] ), .B(\mul_b0/fa1_s1_r[22] ), 
        .Z(n55) );
  HS65_GS_FA1X4 U66 ( .A0(\mul_b0/fa1_s2_r[22] ), .B0(n56), .CI(n55), .CO(n810), .S0(n805) );
  HS65_GS_FA1X4 U67 ( .A0(\mul_b0/fa1_s2_r[23] ), .B0(n58), .CI(n57), .CO(n814), .S0(n809) );
  HS65_GS_FA1X4 U68 ( .A0(\mul_b0/fa1_s2_r[25] ), .B0(n60), .CI(n59), .CO(n822), .S0(n818) );
  HS65_GS_AND2X4 U69 ( .A(\mul_b0/fa1_s1_r[25] ), .B(\mul_b0/fa1_s0_r[25] ), 
        .Z(n62) );
  HS65_GSS_XOR2X3 U70 ( .A(\mul_b0/fa1_s0_r[26] ), .B(\mul_b0/fa1_s1_r[26] ), 
        .Z(n61) );
  HS65_GS_FA1X4 U71 ( .A0(\mul_b0/fa1_s2_r[26] ), .B0(n62), .CI(n61), .CO(n826), .S0(n821) );
  HS65_GS_AND2X4 U72 ( .A(\mul_b0/fa1_s1_r[26] ), .B(\mul_b0/fa1_s0_r[26] ), 
        .Z(n64) );
  HS65_GSS_XOR2X3 U73 ( .A(\mul_b0/fa1_s0_r[27] ), .B(\mul_b0/fa1_s1_r[27] ), 
        .Z(n63) );
  HS65_GS_FA1X4 U74 ( .A0(\mul_b0/fa1_s2_r[27] ), .B0(n64), .CI(n63), .CO(n830), .S0(n825) );
  HS65_GS_FA1X4 U75 ( .A0(\mul_b0/fa1_s2_r[28] ), .B0(n66), .CI(n65), .CO(n534), .S0(n829) );
  HS65_GS_IVX2 U76 ( .A(n67), .Z(n537) );
  HS65_GSS_XOR2X3 U77 ( .A(\mul_b0/fa1_s0_r[31] ), .B(\mul_b0/fa1_s1_r[31] ), 
        .Z(n74) );
  HS65_GS_AND2X4 U78 ( .A(\mul_b0/fa1_s1_r[30] ), .B(\mul_b0/fa1_s0_r[30] ), 
        .Z(n73) );
  HS65_GS_FA1X4 U79 ( .A0(\mul_b0/fa1_s2_r[30] ), .B0(n69), .CI(n68), .CO(n70), 
        .S0(n530) );
  HS65_GS_NAND2X2 U80 ( .A(n71), .B(n70), .Z(n72) );
  HS65_GS_OAI21X2 U81 ( .A(n71), .B(n70), .C(n72), .Z(n536) );
  HS65_GS_NOR2X2 U82 ( .A(n537), .B(n536), .Z(n535) );
  HS65_GS_IVX2 U83 ( .A(n72), .Z(n77) );
  HS65_GSS_XOR2X3 U84 ( .A(\mul_b0/fa1_s0_r[32] ), .B(\mul_b0/fa1_s1_r[32] ), 
        .Z(n80) );
  HS65_GS_AND2X4 U85 ( .A(\mul_b0/fa1_s1_r[31] ), .B(\mul_b0/fa1_s0_r[31] ), 
        .Z(n79) );
  HS65_GS_FA1X4 U86 ( .A0(\mul_b0/fa1_s2_r[31] ), .B0(n74), .CI(n73), .CO(n75), 
        .S0(n71) );
  HS65_GS_FA1X4 U87 ( .A0(n77), .B0(n76), .CI(n75), .CO(n78), .S0(n528) );
  HS65_GS_AOI12X2 U88 ( .A(n535), .B(n528), .C(n78), .Z(n85) );
  HS65_GS_AND2X4 U89 ( .A(\mul_b0/fa1_s1_r[32] ), .B(\mul_b0/fa1_s0_r[32] ), 
        .Z(n82) );
  HS65_GS_FA1X4 U90 ( .A0(\mul_b0/fa1_s2_r[32] ), .B0(n80), .CI(n79), .CO(n81), 
        .S0(n76) );
  HS65_GSS_XOR3X2 U91 ( .A(n82), .B(n81), .C(\mul_b0/fa1_s2_r[33] ), .Z(n83)
         );
  HS65_GSS_XOR3X2 U92 ( .A(\mul_b0/fa1_s0_r[33] ), .B(\mul_b0/fa1_s1_r[33] ), 
        .C(n83), .Z(n84) );
  HS65_GSS_XNOR2X3 U93 ( .A(n85), .B(n84), .Z(\mul_b0/result_sat[15] ) );
  HS65_GS_AND2X4 U94 ( .A(\mul_b1/fa1_c1_r[28] ), .B(\mul_b1/fa1_s2_r[29] ), 
        .Z(n262) );
  HS65_GSS_XOR2X3 U95 ( .A(\mul_b1/fa1_c1_r[28] ), .B(\mul_b1/fa1_s2_r[29] ), 
        .Z(n88) );
  HS65_GSS_XOR2X3 U96 ( .A(\mul_b1/fa1_s0_r[29] ), .B(\mul_b1/fa1_c0_r[28] ), 
        .Z(n87) );
  HS65_GS_AND2X4 U97 ( .A(\mul_b1/fa1_s0_r[28] ), .B(\mul_b1/fa1_c0_r[27] ), 
        .Z(n86) );
  HS65_GS_AND2X4 U98 ( .A(\mul_b1/fa1_s0_r[29] ), .B(\mul_b1/fa1_c0_r[28] ), 
        .Z(n265) );
  HS65_GSS_XOR2X3 U99 ( .A(\mul_b1/fa1_c1_r[29] ), .B(\mul_b1/fa1_s2_r[30] ), 
        .Z(n264) );
  HS65_GSS_XOR2X3 U100 ( .A(\mul_b1/fa1_s0_r[30] ), .B(\mul_b1/fa1_c0_r[29] ), 
        .Z(n263) );
  HS65_GS_AND2X4 U101 ( .A(\mul_b1/fa1_c1_r[27] ), .B(\mul_b1/fa1_s2_r[28] ), 
        .Z(n259) );
  HS65_GSS_XOR2X3 U102 ( .A(\mul_b1/fa1_s0_r[28] ), .B(\mul_b1/fa1_c0_r[27] ), 
        .Z(n91) );
  HS65_GSS_XOR2X3 U103 ( .A(\mul_b1/fa1_c1_r[27] ), .B(\mul_b1/fa1_s2_r[28] ), 
        .Z(n90) );
  HS65_GS_AND2X4 U104 ( .A(\mul_b1/fa1_s0_r[27] ), .B(\mul_b1/fa1_c0_r[26] ), 
        .Z(n89) );
  HS65_GS_FA1X4 U105 ( .A0(n88), .B0(n87), .CI(n86), .CO(n261), .S0(n257) );
  HS65_GS_AND2X4 U106 ( .A(\mul_b1/fa1_c1_r[26] ), .B(\mul_b1/fa1_s2_r[27] ), 
        .Z(n256) );
  HS65_GSS_XOR2X3 U107 ( .A(\mul_b1/fa1_s0_r[27] ), .B(\mul_b1/fa1_c0_r[26] ), 
        .Z(n94) );
  HS65_GSS_XOR2X3 U108 ( .A(\mul_b1/fa1_c1_r[26] ), .B(\mul_b1/fa1_s2_r[27] ), 
        .Z(n93) );
  HS65_GS_AND2X4 U109 ( .A(\mul_b1/fa1_s0_r[26] ), .B(\mul_b1/fa1_c0_r[25] ), 
        .Z(n92) );
  HS65_GS_FA1X4 U110 ( .A0(n91), .B0(n90), .CI(n89), .CO(n258), .S0(n254) );
  HS65_GS_AND2X4 U111 ( .A(\mul_b1/fa1_c1_r[25] ), .B(\mul_b1/fa1_s2_r[26] ), 
        .Z(n97) );
  HS65_GSS_XOR2X3 U112 ( .A(\mul_b1/fa1_s0_r[26] ), .B(\mul_b1/fa1_c0_r[25] ), 
        .Z(n250) );
  HS65_GSS_XOR2X3 U113 ( .A(\mul_b1/fa1_c1_r[25] ), .B(\mul_b1/fa1_s2_r[26] ), 
        .Z(n249) );
  HS65_GS_AND2X4 U114 ( .A(\mul_b1/fa1_s0_r[25] ), .B(\mul_b1/fa1_c0_r[24] ), 
        .Z(n248) );
  HS65_GS_FA1X4 U115 ( .A0(n94), .B0(n93), .CI(n92), .CO(n255), .S0(n95) );
  HS65_GS_FA1X4 U116 ( .A0(n97), .B0(n96), .CI(n95), .CO(n931), .S0(n928) );
  HS65_GSS_XOR2X3 U117 ( .A(\mul_b1/fa1_c1_r[22] ), .B(\mul_b1/fa1_s2_r[23] ), 
        .Z(n104) );
  HS65_GSS_XOR2X3 U118 ( .A(\mul_b1/fa1_s0_r[23] ), .B(\mul_b1/fa1_c0_r[22] ), 
        .Z(n103) );
  HS65_GS_AOI12X2 U119 ( .A(\mul_b1/fa1_s2_r[23] ), .B(\mul_b1/fa1_c1_r[22] ), 
        .C(n100), .Z(n101) );
  HS65_GSS_XOR2X3 U120 ( .A(\mul_b1/fa1_s0_r[24] ), .B(\mul_b1/fa1_c0_r[23] ), 
        .Z(n241) );
  HS65_GSS_XOR2X3 U121 ( .A(\mul_b1/fa1_c1_r[23] ), .B(\mul_b1/fa1_s2_r[24] ), 
        .Z(n240) );
  HS65_GS_AND2X4 U122 ( .A(\mul_b1/fa1_s0_r[23] ), .B(\mul_b1/fa1_c0_r[22] ), 
        .Z(n239) );
  HS65_GS_AND2X4 U123 ( .A(\mul_b1/fa1_c1_r[22] ), .B(\mul_b1/fa1_s2_r[23] ), 
        .Z(n99) );
  HS65_GS_NAND3X2 U124 ( .A(n103), .B(n102), .C(n99), .Z(n98) );
  HS65_GS_OAI21X2 U125 ( .A(n100), .B(n99), .C(n98), .Z(n237) );
  HS65_GS_NOR2X2 U126 ( .A(n238), .B(n237), .Z(n236) );
  HS65_GS_NOR2X2 U127 ( .A(n101), .B(n236), .Z(n922) );
  HS65_GS_AND2X4 U128 ( .A(\mul_b1/fa1_c1_r[21] ), .B(\mul_b1/fa1_s2_r[22] ), 
        .Z(n235) );
  HS65_GSS_XOR2X3 U129 ( .A(\mul_b1/fa1_c1_r[21] ), .B(\mul_b1/fa1_s2_r[22] ), 
        .Z(n108) );
  HS65_GS_FA1X4 U130 ( .A0(\mul_b1/fa1_s0_r[22] ), .B0(\mul_b1/fa1_s1_r[22] ), 
        .CI(\mul_b1/fa1_c0_r[21] ), .CO(n102), .S0(n106) );
  HS65_GS_FA1X4 U131 ( .A0(n104), .B0(n103), .CI(n102), .CO(n100), .S0(n233)
         );
  HS65_GS_FA1X4 U132 ( .A0(\mul_b1/fa1_s0_r[21] ), .B0(\mul_b1/fa1_s1_r[21] ), 
        .CI(\mul_b1/fa1_c0_r[20] ), .CO(n107), .S0(n119) );
  HS65_GS_NAND2X2 U133 ( .A(n120), .B(n119), .Z(n118) );
  HS65_GS_IVX2 U134 ( .A(n118), .Z(n110) );
  HS65_GS_FA1X4 U135 ( .A0(\mul_b1/fa1_s2_r[21] ), .B0(\mul_b1/fa1_c1_r[20] ), 
        .CI(n105), .CO(n111), .S0(n120) );
  HS65_GS_NOR2X2 U136 ( .A(n110), .B(n111), .Z(n112) );
  HS65_GS_FA1X4 U137 ( .A0(n108), .B0(n107), .CI(n106), .CO(n234), .S0(n232)
         );
  HS65_GS_NAND3X2 U138 ( .A(\mul_b1/fa1_s2_r[21] ), .B(\mul_b1/fa1_c1_r[20] ), 
        .C(n110), .Z(n109) );
  HS65_GS_OAI21X2 U139 ( .A(n111), .B(n110), .C(n109), .Z(n231) );
  HS65_GS_NOR2X2 U140 ( .A(n232), .B(n231), .Z(n230) );
  HS65_GS_NOR2X2 U141 ( .A(n112), .B(n230), .Z(n914) );
  HS65_GS_NAND2X2 U142 ( .A(\mul_b1/fa1_c1_r[19] ), .B(\mul_b1/fa1_s2_r[20] ), 
        .Z(n113) );
  HS65_GS_IVX2 U143 ( .A(n113), .Z(n116) );
  HS65_GS_FA1X4 U144 ( .A0(\mul_b1/fa1_s0_r[20] ), .B0(\mul_b1/fa1_s1_r[20] ), 
        .CI(\mul_b1/fa1_c0_r[19] ), .CO(n105), .S0(n126) );
  HS65_GS_OA12X4 U145 ( .A(\mul_b1/fa1_c1_r[19] ), .B(\mul_b1/fa1_s2_r[20] ), 
        .C(n113), .Z(n114) );
  HS65_GS_AND2X4 U146 ( .A(n117), .B(n114), .Z(n127) );
  HS65_GS_NOR2X2 U147 ( .A(n117), .B(n114), .Z(n125) );
  HS65_GS_NOR2AX3 U148 ( .A(n126), .B(n125), .Z(n115) );
  HS65_GS_NOR3X1 U149 ( .A(n116), .B(n127), .C(n115), .Z(n121) );
  HS65_GS_AOI13X2 U150 ( .A(n117), .B(n116), .C(n126), .D(n121), .Z(n229) );
  HS65_GS_OAI21X2 U151 ( .A(n120), .B(n119), .C(n118), .Z(n228) );
  HS65_GS_NAND2X2 U152 ( .A(n229), .B(n228), .Z(n227) );
  HS65_GS_NOR2AX3 U153 ( .A(n227), .B(n121), .Z(n910) );
  HS65_GS_IVX2 U154 ( .A(n122), .Z(n136) );
  HS65_GS_NAND2X2 U155 ( .A(\mul_b1/fa1_c1_r[18] ), .B(\mul_b1/fa1_s2_r[19] ), 
        .Z(n128) );
  HS65_GS_OAI21X2 U156 ( .A(\mul_b1/fa1_c1_r[18] ), .B(\mul_b1/fa1_s2_r[19] ), 
        .C(n128), .Z(n123) );
  HS65_GS_IVX2 U157 ( .A(n123), .Z(n134) );
  HS65_GS_FA1X4 U158 ( .A0(\mul_b1/fa1_s0_r[19] ), .B0(\mul_b1/fa1_s1_r[19] ), 
        .CI(\mul_b1/fa1_c0_r[18] ), .CO(n117), .S0(n135) );
  HS65_GS_OAI21X2 U159 ( .A(n122), .B(n134), .C(n135), .Z(n129) );
  HS65_GS_OAI112X1 U160 ( .A(n136), .B(n123), .C(n128), .D(n129), .Z(n130) );
  HS65_GS_OAI21X2 U161 ( .A(n127), .B(n125), .C(n126), .Z(n124) );
  HS65_GS_OAI13X1 U162 ( .A(n127), .B(n126), .C(n125), .D(n124), .Z(n226) );
  HS65_GS_OAI21X2 U163 ( .A(n129), .B(n128), .C(n130), .Z(n225) );
  HS65_GS_NOR2X2 U164 ( .A(n226), .B(n225), .Z(n224) );
  HS65_GS_NOR2AX3 U165 ( .A(n130), .B(n224), .Z(n906) );
  HS65_GS_FA1X4 U166 ( .A0(\mul_b1/fa1_s0_r[18] ), .B0(\mul_b1/fa1_s1_r[18] ), 
        .CI(\mul_b1/fa1_c0_r[17] ), .CO(n122), .S0(n143) );
  HS65_GS_NAND2X2 U167 ( .A(n144), .B(n143), .Z(n142) );
  HS65_GS_IVX2 U168 ( .A(n142), .Z(n133) );
  HS65_GS_FA1X4 U169 ( .A0(\mul_b1/fa1_s2_r[18] ), .B0(\mul_b1/fa1_c1_r[17] ), 
        .CI(n131), .CO(n132), .S0(n144) );
  HS65_GS_AOI12X2 U170 ( .A(n143), .B(n144), .C(n132), .Z(n137) );
  HS65_GS_AOI13X2 U171 ( .A(n133), .B(\mul_b1/fa1_c1_r[17] ), .C(
        \mul_b1/fa1_s2_r[18] ), .D(n137), .Z(n139) );
  HS65_GSS_XOR3X2 U172 ( .A(n136), .B(n135), .C(n134), .Z(n138) );
  HS65_GS_AOI12X2 U173 ( .A(n139), .B(n138), .C(n137), .Z(n902) );
  HS65_GSS_XOR2X3 U174 ( .A(n139), .B(n138), .Z(n569) );
  HS65_GS_FA1X4 U175 ( .A0(\mul_b1/fa1_s0_r[17] ), .B0(\mul_b1/fa1_s1_r[17] ), 
        .CI(\mul_b1/fa1_c0_r[16] ), .CO(n131), .S0(n151) );
  HS65_GS_NAND2X2 U176 ( .A(n152), .B(n151), .Z(n150) );
  HS65_GS_IVX2 U177 ( .A(n150), .Z(n146) );
  HS65_GS_FA1X4 U178 ( .A0(\mul_b1/fa1_s2_r[17] ), .B0(\mul_b1/fa1_c1_r[16] ), 
        .CI(n140), .CO(n145), .S0(n152) );
  HS65_GS_AOI12X2 U179 ( .A(n151), .B(n152), .C(n145), .Z(n141) );
  HS65_GS_AOI13X2 U180 ( .A(n146), .B(\mul_b1/fa1_c1_r[16] ), .C(
        \mul_b1/fa1_s2_r[17] ), .D(n141), .Z(n156) );
  HS65_GS_OAI21X2 U181 ( .A(n144), .B(n143), .C(n142), .Z(n155) );
  HS65_GS_NAND2X2 U182 ( .A(n156), .B(n155), .Z(n154) );
  HS65_GS_OAI21X2 U183 ( .A(n146), .B(n145), .C(n154), .Z(n547) );
  HS65_GS_FA1X4 U184 ( .A0(\mul_b1/fa1_s0_r[16] ), .B0(\mul_b1/fa1_s1_r[16] ), 
        .CI(\mul_b1/fa1_c0_r[15] ), .CO(n140), .S0(n161) );
  HS65_GS_NAND2X2 U185 ( .A(n162), .B(n161), .Z(n160) );
  HS65_GS_IVX2 U186 ( .A(n160), .Z(n149) );
  HS65_GS_FA1X4 U187 ( .A0(\mul_b1/fa1_s2_r[16] ), .B0(\mul_b1/fa1_c1_r[15] ), 
        .CI(n147), .CO(n148), .S0(n162) );
  HS65_GS_AOI12X2 U188 ( .A(n161), .B(n162), .C(n148), .Z(n153) );
  HS65_GS_AOI13X2 U189 ( .A(n149), .B(\mul_b1/fa1_s2_r[16] ), .C(
        \mul_b1/fa1_c1_r[15] ), .D(n153), .Z(n222) );
  HS65_GS_OAI21X2 U190 ( .A(n152), .B(n151), .C(n150), .Z(n221) );
  HS65_GS_NAND2X2 U191 ( .A(n222), .B(n221), .Z(n220) );
  HS65_GS_NOR2AX3 U192 ( .A(n220), .B(n153), .Z(n898) );
  HS65_GS_OAI21X2 U193 ( .A(n156), .B(n155), .C(n154), .Z(n897) );
  HS65_GS_FA1X4 U194 ( .A0(\mul_b1/fa1_s0_r[15] ), .B0(\mul_b1/fa1_s1_r[15] ), 
        .CI(\mul_b1/fa1_c0_r[14] ), .CO(n147), .S0(n157) );
  HS65_GS_AND2X4 U195 ( .A(n166), .B(n165), .Z(n159) );
  HS65_GS_FA1X4 U196 ( .A0(\mul_b1/fa1_s2_r[15] ), .B0(\mul_b1/fa1_c1_r[14] ), 
        .CI(n157), .CO(n158), .S0(n166) );
  HS65_GS_AOI12X2 U197 ( .A(n165), .B(n166), .C(n158), .Z(n218) );
  HS65_GS_AOI13X2 U198 ( .A(n159), .B(\mul_b1/fa1_s2_r[15] ), .C(
        \mul_b1/fa1_c1_r[14] ), .D(n218), .Z(n164) );
  HS65_GS_OAI21X2 U199 ( .A(n162), .B(n161), .C(n160), .Z(n163) );
  HS65_GS_NAND2X2 U200 ( .A(n164), .B(n163), .Z(n219) );
  HS65_GS_OAI21X2 U201 ( .A(n164), .B(n163), .C(n219), .Z(n890) );
  HS65_GS_AND2X4 U202 ( .A(\mul_b1/fa1_c1_r[13] ), .B(\mul_b1/fa1_s2_r[14] ), 
        .Z(n169) );
  HS65_GSS_XOR2X3 U203 ( .A(n166), .B(n165), .Z(n168) );
  HS65_GSS_XOR2X3 U204 ( .A(\mul_b1/fa1_c1_r[13] ), .B(\mul_b1/fa1_s2_r[14] ), 
        .Z(n211) );
  HS65_GS_FA1X4 U205 ( .A0(\mul_b1/fa1_s0_r[14] ), .B0(\mul_b1/fa1_s1_r[14] ), 
        .CI(\mul_b1/fa1_c0_r[13] ), .CO(n165), .S0(n210) );
  HS65_GS_FA1X4 U206 ( .A0(n169), .B0(n168), .CI(n167), .CO(n889), .S0(n886)
         );
  HS65_GS_FA1X4 U207 ( .A0(\mul_b1/fa1_s0_r[13] ), .B0(\mul_b1/fa1_s1_r[13] ), 
        .CI(\mul_b1/fa1_c0_r[12] ), .CO(n209), .S0(n213) );
  HS65_GSS_XOR2X3 U208 ( .A(\mul_b1/fa1_c1_r[12] ), .B(\mul_b1/fa1_s2_r[13] ), 
        .Z(n212) );
  HS65_GS_FA1X4 U209 ( .A0(\mul_b1/fa1_s0_r[12] ), .B0(\mul_b1/fa1_s1_r[12] ), 
        .CI(\mul_b1/fa1_c0_r[11] ), .CO(n214), .S0(n175) );
  HS65_GS_NAND2X2 U210 ( .A(n176), .B(n175), .Z(n174) );
  HS65_GS_IVX2 U211 ( .A(n174), .Z(n172) );
  HS65_GS_FA1X4 U212 ( .A0(\mul_b1/fa1_s2_r[12] ), .B0(\mul_b1/fa1_c1_r[11] ), 
        .CI(n170), .CO(n171), .S0(n176) );
  HS65_GS_AOI12X2 U213 ( .A(n175), .B(n176), .C(n171), .Z(n206) );
  HS65_GS_AOI13X2 U214 ( .A(n172), .B(\mul_b1/fa1_s2_r[12] ), .C(
        \mul_b1/fa1_c1_r[11] ), .D(n206), .Z(n208) );
  HS65_GS_FA1X4 U215 ( .A0(\mul_b1/fa1_s0_r[11] ), .B0(\mul_b1/fa1_s1_r[11] ), 
        .CI(\mul_b1/fa1_c0_r[10] ), .CO(n170), .S0(n177) );
  HS65_GS_IVX2 U216 ( .A(n173), .Z(n202) );
  HS65_GS_OAI21X2 U217 ( .A(n176), .B(n175), .C(n174), .Z(n201) );
  HS65_GS_FA1X4 U218 ( .A0(\mul_b1/fa1_s0_r[10] ), .B0(\mul_b1/fa1_s1_r[10] ), 
        .CI(\mul_b1/fa1_c0_r[9] ), .CO(n178), .S0(n188) );
  HS65_GS_FA1X4 U219 ( .A0(\mul_b1/fa1_c1_r[10] ), .B0(n178), .CI(n177), .CO(
        n173), .S0(n198) );
  HS65_GS_FA1X4 U220 ( .A0(\mul_b1/fa1_s0_r[7] ), .B0(\mul_b1/fa1_s1_r[7] ), 
        .CI(\mul_b1/fa1_c0_r[6] ), .CO(n185), .S0(n183) );
  HS65_GS_OAI112X1 U221 ( .A(\mul_b1/fa1_c0_r[4] ), .B(\mul_b1/fa1_s0_r[5] ), 
        .C(\mul_b1/fa1_c0_r[3] ), .D(\mul_b1/fa1_s0_r[4] ), .Z(n180) );
  HS65_GS_NAND2X2 U222 ( .A(\mul_b1/fa1_s0_r[5] ), .B(\mul_b1/fa1_c0_r[4] ), 
        .Z(n179) );
  HS65_GS_NAND2X2 U223 ( .A(n180), .B(n179), .Z(n181) );
  HS65_GS_PAOI2X1 U224 ( .A(\mul_b1/fa1_c0_r[5] ), .B(\mul_b1/fa1_s0_r[6] ), 
        .P(n181), .Z(n182) );
  HS65_GS_NOR2AX3 U225 ( .A(n183), .B(n182), .Z(n184) );
  HS65_GS_PAOI2X1 U226 ( .A(n186), .B(n185), .P(n184), .Z(n196) );
  HS65_GS_FA1X4 U227 ( .A0(\mul_b1/fa1_s0_r[8] ), .B0(\mul_b1/fa1_s1_r[8] ), 
        .CI(\mul_b1/fa1_c0_r[7] ), .CO(n190), .S0(n186) );
  HS65_GS_FA1X4 U228 ( .A0(\mul_b1/fa1_s0_r[9] ), .B0(\mul_b1/fa1_s1_r[9] ), 
        .CI(\mul_b1/fa1_c0_r[8] ), .CO(n187), .S0(n189) );
  HS65_GS_FA1X4 U229 ( .A0(\mul_b1/fa1_c1_r[9] ), .B0(n188), .CI(n187), .CO(
        n199), .S0(n192) );
  HS65_GS_FA1X4 U230 ( .A0(\mul_b1/fa1_c1_r[8] ), .B0(n190), .CI(n189), .CO(
        n193), .S0(n191) );
  HS65_GS_OAI21X2 U231 ( .A(n193), .B(n192), .C(n191), .Z(n195) );
  HS65_GS_NAND2X2 U232 ( .A(n193), .B(n192), .Z(n194) );
  HS65_GS_OAI21X2 U233 ( .A(n196), .B(n195), .C(n194), .Z(n197) );
  HS65_GS_PAOI2X1 U234 ( .A(n199), .B(n198), .P(n197), .Z(n200) );
  HS65_GS_PAOI2X1 U235 ( .A(n202), .B(n201), .P(n200), .Z(n203) );
  HS65_GS_OAI21X2 U236 ( .A(n205), .B(n208), .C(n203), .Z(n204) );
  HS65_GS_AOI12X2 U237 ( .A(n205), .B(n208), .C(n204), .Z(n882) );
  HS65_GS_IVX2 U238 ( .A(n205), .Z(n207) );
  HS65_GS_AOI12X2 U239 ( .A(n208), .B(n207), .C(n206), .Z(n881) );
  HS65_GS_AND2X4 U240 ( .A(\mul_b1/fa1_c1_r[12] ), .B(\mul_b1/fa1_s2_r[13] ), 
        .Z(n217) );
  HS65_GS_FA1X4 U241 ( .A0(n211), .B0(n210), .CI(n209), .CO(n167), .S0(n216)
         );
  HS65_GS_FA1X4 U242 ( .A0(n214), .B0(n213), .CI(n212), .CO(n215), .S0(n205)
         );
  HS65_GS_FA1X4 U243 ( .A0(n217), .B0(n216), .CI(n215), .CO(n884), .S0(n880)
         );
  HS65_GS_NOR2AX3 U244 ( .A(n219), .B(n218), .Z(n893) );
  HS65_GS_OAI21X2 U245 ( .A(n222), .B(n221), .C(n220), .Z(n892) );
  HS65_GS_IVX2 U246 ( .A(n223), .Z(n548) );
  HS65_GS_PAOI2X1 U247 ( .A(n569), .B(n547), .P(n548), .Z(n901) );
  HS65_GS_AO12X4 U248 ( .A(n226), .B(n225), .C(n224), .Z(n900) );
  HS65_GS_OAI21X2 U249 ( .A(n229), .B(n228), .C(n227), .Z(n904) );
  HS65_GS_AO12X4 U250 ( .A(n232), .B(n231), .C(n230), .Z(n908) );
  HS65_GS_FA1X4 U251 ( .A0(n235), .B0(n234), .CI(n233), .CO(n918), .S0(n912)
         );
  HS65_GS_AO12X4 U252 ( .A(n238), .B(n237), .C(n236), .Z(n916) );
  HS65_GS_AND2X4 U253 ( .A(\mul_b1/fa1_c1_r[23] ), .B(\mul_b1/fa1_s2_r[24] ), 
        .Z(n244) );
  HS65_GS_FA1X4 U254 ( .A0(n241), .B0(n240), .CI(n239), .CO(n243), .S0(n238)
         );
  HS65_GSS_XOR2X3 U255 ( .A(\mul_b1/fa1_s0_r[25] ), .B(\mul_b1/fa1_c0_r[24] ), 
        .Z(n247) );
  HS65_GSS_XOR2X3 U256 ( .A(\mul_b1/fa1_c1_r[24] ), .B(\mul_b1/fa1_s2_r[25] ), 
        .Z(n246) );
  HS65_GS_AND2X4 U257 ( .A(\mul_b1/fa1_s0_r[24] ), .B(\mul_b1/fa1_c0_r[23] ), 
        .Z(n245) );
  HS65_GS_FA1X4 U258 ( .A0(n244), .B0(n243), .CI(n242), .CO(n1033), .S0(n920)
         );
  HS65_GS_AND2X4 U259 ( .A(\mul_b1/fa1_c1_r[24] ), .B(\mul_b1/fa1_s2_r[25] ), 
        .Z(n253) );
  HS65_GS_FA1X4 U260 ( .A0(n247), .B0(n246), .CI(n245), .CO(n252), .S0(n242)
         );
  HS65_GS_FA1X4 U261 ( .A0(n250), .B0(n249), .CI(n248), .CO(n96), .S0(n251) );
  HS65_GS_PAO2X4 U262 ( .A(n1032), .B(n1033), .P(n1035), .Z(n924) );
  HS65_GS_FA1X4 U263 ( .A0(n253), .B0(n252), .CI(n251), .CO(n925), .S0(n1035)
         );
  HS65_GS_PAO2X4 U264 ( .A(n928), .B(n924), .P(n925), .Z(n930) );
  HS65_GS_FA1X4 U265 ( .A0(n256), .B0(n255), .CI(n254), .CO(n558), .S0(n929)
         );
  HS65_GS_FA1X4 U266 ( .A0(n259), .B0(n258), .CI(n257), .CO(n561), .S0(n556)
         );
  HS65_GS_FA1X4 U267 ( .A0(n262), .B0(n261), .CI(n260), .CO(n555), .S0(n559)
         );
  HS65_GS_FA1X4 U268 ( .A0(n265), .B0(n264), .CI(n263), .CO(n271), .S0(n260)
         );
  HS65_GS_AND2X4 U269 ( .A(\mul_b1/fa1_c1_r[29] ), .B(\mul_b1/fa1_s2_r[30] ), 
        .Z(n270) );
  HS65_GS_AND2X4 U270 ( .A(\mul_b1/fa1_s0_r[30] ), .B(\mul_b1/fa1_c0_r[29] ), 
        .Z(n268) );
  HS65_GSS_XOR2X3 U271 ( .A(\mul_b1/fa1_c1_r[30] ), .B(\mul_b1/fa1_s2_r[31] ), 
        .Z(n267) );
  HS65_GSS_XOR2X3 U272 ( .A(\mul_b1/fa1_s0_r[31] ), .B(\mul_b1/fa1_c0_r[30] ), 
        .Z(n266) );
  HS65_GS_AND2X4 U273 ( .A(\mul_b1/fa1_c1_r[30] ), .B(\mul_b1/fa1_s2_r[31] ), 
        .Z(n274) );
  HS65_GS_AND2X4 U274 ( .A(\mul_b1/fa1_s0_r[31] ), .B(\mul_b1/fa1_c0_r[30] ), 
        .Z(n277) );
  HS65_GS_NAND2X2 U275 ( .A(\mul_b1/fa1_c1_r[31] ), .B(\mul_b1/fa1_s2_r[32] ), 
        .Z(n278) );
  HS65_GS_OA12X4 U276 ( .A(\mul_b1/fa1_c1_r[31] ), .B(\mul_b1/fa1_s2_r[32] ), 
        .C(n278), .Z(n276) );
  HS65_GS_NAND2X2 U277 ( .A(\mul_b1/fa1_s0_r[32] ), .B(\mul_b1/fa1_c0_r[31] ), 
        .Z(n280) );
  HS65_GS_OA12X4 U278 ( .A(\mul_b1/fa1_s0_r[32] ), .B(\mul_b1/fa1_c0_r[31] ), 
        .C(n280), .Z(n275) );
  HS65_GS_FA1X4 U279 ( .A0(n268), .B0(n267), .CI(n266), .CO(n272), .S0(n269)
         );
  HS65_GS_FA1X4 U280 ( .A0(n271), .B0(n270), .CI(n269), .CO(n549), .S0(n553)
         );
  HS65_GS_FA1X4 U281 ( .A0(n274), .B0(n273), .CI(n272), .CO(n283), .S0(n550)
         );
  HS65_GS_FA1X4 U282 ( .A0(n277), .B0(n276), .CI(n275), .CO(n281), .S0(n273)
         );
  HS65_GSS_XOR3X2 U283 ( .A(\mul_b1/fa1_s2_r[33] ), .B(\mul_b1/fa1_s0_r[33] ), 
        .C(n278), .Z(n279) );
  HS65_GSS_XOR3X2 U284 ( .A(n281), .B(n280), .C(n279), .Z(n282) );
  HS65_GSS_XOR3X2 U285 ( .A(n284), .B(n283), .C(n282), .Z(n285) );
  HS65_GSS_XOR3X2 U286 ( .A(\mul_b1/fa1_c0_r[32] ), .B(\mul_b1/fa1_c1_r[32] ), 
        .C(n285), .Z(\mul_b1/result_sat[15] ) );
  HS65_GS_AND2X4 U287 ( .A(\mul_a1/fa1_c1_r[31] ), .B(\mul_a1/fa1_s2_r[32] ), 
        .Z(n450) );
  HS65_GS_FA1X4 U288 ( .A0(\mul_a1/fa1_c1_r[27] ), .B0(\mul_a1/fa1_c2_r[27] ), 
        .CI(\mul_a1/fa1_s2_r[28] ), .CO(n420), .S0(n288) );
  HS65_GSS_XOR2X3 U289 ( .A(\mul_a1/fa1_s0_r[28] ), .B(\mul_a1/fa1_s1_r[28] ), 
        .Z(n287) );
  HS65_GS_AND2X4 U290 ( .A(\mul_a1/fa1_s0_r[27] ), .B(\mul_a1/fa1_s1_r[27] ), 
        .Z(n286) );
  HS65_GS_AND2X4 U291 ( .A(\mul_a1/fa1_s0_r[28] ), .B(\mul_a1/fa1_s1_r[28] ), 
        .Z(n423) );
  HS65_GSS_XOR2X3 U292 ( .A(\mul_a1/fa1_s0_r[29] ), .B(\mul_a1/fa1_s1_r[29] ), 
        .Z(n421) );
  HS65_GS_FA1X4 U293 ( .A0(\mul_a1/fa1_c1_r[26] ), .B0(\mul_a1/fa1_c2_r[26] ), 
        .CI(\mul_a1/fa1_s2_r[27] ), .CO(n417), .S0(n291) );
  HS65_GSS_XOR2X3 U294 ( .A(\mul_a1/fa1_s0_r[27] ), .B(\mul_a1/fa1_s1_r[27] ), 
        .Z(n290) );
  HS65_GS_AND2X4 U295 ( .A(\mul_a1/fa1_s0_r[26] ), .B(\mul_a1/fa1_s1_r[26] ), 
        .Z(n289) );
  HS65_GS_FA1X4 U296 ( .A0(n288), .B0(n287), .CI(n286), .CO(n419), .S0(n415)
         );
  HS65_GS_FA1X4 U297 ( .A0(\mul_a1/fa1_c1_r[25] ), .B0(\mul_a1/fa1_c2_r[25] ), 
        .CI(\mul_a1/fa1_s2_r[26] ), .CO(n414), .S0(n294) );
  HS65_GSS_XOR2X3 U298 ( .A(\mul_a1/fa1_s0_r[26] ), .B(\mul_a1/fa1_s1_r[26] ), 
        .Z(n293) );
  HS65_GS_AND2X4 U299 ( .A(\mul_a1/fa1_s0_r[25] ), .B(\mul_a1/fa1_s1_r[25] ), 
        .Z(n292) );
  HS65_GS_FA1X4 U300 ( .A0(n291), .B0(n290), .CI(n289), .CO(n416), .S0(n412)
         );
  HS65_GS_FA1X4 U301 ( .A0(\mul_a1/fa1_c1_r[24] ), .B0(\mul_a1/fa1_c2_r[24] ), 
        .CI(\mul_a1/fa1_s2_r[25] ), .CO(n411), .S0(n297) );
  HS65_GSS_XOR2X3 U302 ( .A(\mul_a1/fa1_s0_r[25] ), .B(\mul_a1/fa1_s1_r[25] ), 
        .Z(n296) );
  HS65_GS_AND2X4 U303 ( .A(\mul_a1/fa1_s0_r[24] ), .B(\mul_a1/fa1_s1_r[24] ), 
        .Z(n295) );
  HS65_GS_FA1X4 U304 ( .A0(n294), .B0(n293), .CI(n292), .CO(n413), .S0(n409)
         );
  HS65_GS_FA1X4 U305 ( .A0(\mul_a1/fa1_c1_r[23] ), .B0(\mul_a1/fa1_c2_r[23] ), 
        .CI(\mul_a1/fa1_s2_r[24] ), .CO(n408), .S0(n300) );
  HS65_GSS_XOR2X3 U306 ( .A(\mul_a1/fa1_s0_r[24] ), .B(\mul_a1/fa1_s1_r[24] ), 
        .Z(n299) );
  HS65_GS_AND2X4 U307 ( .A(\mul_a1/fa1_s0_r[23] ), .B(\mul_a1/fa1_s1_r[23] ), 
        .Z(n298) );
  HS65_GS_FA1X4 U308 ( .A0(n297), .B0(n296), .CI(n295), .CO(n410), .S0(n406)
         );
  HS65_GS_FA1X4 U309 ( .A0(\mul_a1/fa1_c1_r[22] ), .B0(\mul_a1/fa1_c2_r[22] ), 
        .CI(\mul_a1/fa1_s2_r[23] ), .CO(n405), .S0(n303) );
  HS65_GSS_XOR2X3 U310 ( .A(\mul_a1/fa1_s0_r[23] ), .B(\mul_a1/fa1_s1_r[23] ), 
        .Z(n302) );
  HS65_GS_AND2X4 U311 ( .A(\mul_a1/fa1_s0_r[22] ), .B(\mul_a1/fa1_s1_r[22] ), 
        .Z(n301) );
  HS65_GS_FA1X4 U312 ( .A0(n300), .B0(n299), .CI(n298), .CO(n407), .S0(n403)
         );
  HS65_GS_FA1X4 U313 ( .A0(\mul_a1/fa1_c1_r[21] ), .B0(\mul_a1/fa1_c2_r[21] ), 
        .CI(\mul_a1/fa1_s2_r[22] ), .CO(n402), .S0(n306) );
  HS65_GSS_XOR2X3 U314 ( .A(\mul_a1/fa1_s0_r[22] ), .B(\mul_a1/fa1_s1_r[22] ), 
        .Z(n305) );
  HS65_GS_AND2X4 U315 ( .A(\mul_a1/fa1_s0_r[21] ), .B(\mul_a1/fa1_s1_r[21] ), 
        .Z(n304) );
  HS65_GS_FA1X4 U316 ( .A0(n303), .B0(n302), .CI(n301), .CO(n404), .S0(n400)
         );
  HS65_GS_FA1X4 U317 ( .A0(\mul_a1/fa1_c1_r[20] ), .B0(\mul_a1/fa1_c2_r[20] ), 
        .CI(\mul_a1/fa1_s2_r[21] ), .CO(n399), .S0(n309) );
  HS65_GSS_XOR2X3 U318 ( .A(\mul_a1/fa1_s0_r[21] ), .B(\mul_a1/fa1_s1_r[21] ), 
        .Z(n308) );
  HS65_GS_AND2X4 U319 ( .A(\mul_a1/fa1_s0_r[20] ), .B(\mul_a1/fa1_s1_r[20] ), 
        .Z(n307) );
  HS65_GS_FA1X4 U320 ( .A0(n306), .B0(n305), .CI(n304), .CO(n401), .S0(n397)
         );
  HS65_GS_FA1X4 U321 ( .A0(\mul_a1/fa1_c1_r[19] ), .B0(\mul_a1/fa1_c2_r[19] ), 
        .CI(\mul_a1/fa1_s2_r[20] ), .CO(n396), .S0(n312) );
  HS65_GSS_XOR2X3 U322 ( .A(\mul_a1/fa1_s0_r[20] ), .B(\mul_a1/fa1_s1_r[20] ), 
        .Z(n311) );
  HS65_GS_AND2X4 U323 ( .A(\mul_a1/fa1_s0_r[19] ), .B(\mul_a1/fa1_s1_r[19] ), 
        .Z(n310) );
  HS65_GS_FA1X4 U324 ( .A0(n309), .B0(n308), .CI(n307), .CO(n398), .S0(n394)
         );
  HS65_GS_FA1X4 U325 ( .A0(\mul_a1/fa1_c1_r[18] ), .B0(\mul_a1/fa1_c2_r[18] ), 
        .CI(\mul_a1/fa1_s2_r[19] ), .CO(n393), .S0(n315) );
  HS65_GSS_XOR2X3 U326 ( .A(\mul_a1/fa1_s0_r[19] ), .B(\mul_a1/fa1_s1_r[19] ), 
        .Z(n314) );
  HS65_GS_AND2X4 U327 ( .A(\mul_a1/fa1_s0_r[18] ), .B(\mul_a1/fa1_s1_r[18] ), 
        .Z(n313) );
  HS65_GS_FA1X4 U328 ( .A0(n312), .B0(n311), .CI(n310), .CO(n395), .S0(n391)
         );
  HS65_GS_FA1X4 U329 ( .A0(\mul_a1/fa1_c1_r[17] ), .B0(\mul_a1/fa1_c2_r[17] ), 
        .CI(\mul_a1/fa1_s2_r[18] ), .CO(n390), .S0(n318) );
  HS65_GSS_XOR2X3 U330 ( .A(\mul_a1/fa1_s0_r[18] ), .B(\mul_a1/fa1_s1_r[18] ), 
        .Z(n317) );
  HS65_GS_AND2X4 U331 ( .A(\mul_a1/fa1_s0_r[17] ), .B(\mul_a1/fa1_s1_r[17] ), 
        .Z(n316) );
  HS65_GS_FA1X4 U332 ( .A0(n315), .B0(n314), .CI(n313), .CO(n392), .S0(n388)
         );
  HS65_GS_FA1X4 U333 ( .A0(\mul_a1/fa1_c1_r[16] ), .B0(\mul_a1/fa1_c2_r[16] ), 
        .CI(\mul_a1/fa1_s2_r[17] ), .CO(n387), .S0(n376) );
  HS65_GSS_XOR2X3 U334 ( .A(\mul_a1/fa1_s0_r[17] ), .B(\mul_a1/fa1_s1_r[17] ), 
        .Z(n375) );
  HS65_GS_AND2X4 U335 ( .A(\mul_a1/fa1_s0_r[16] ), .B(\mul_a1/fa1_s1_r[16] ), 
        .Z(n374) );
  HS65_GS_FA1X4 U336 ( .A0(n318), .B0(n317), .CI(n316), .CO(n389), .S0(n385)
         );
  HS65_GS_FA1X4 U337 ( .A0(\mul_a1/fa1_c1_r[14] ), .B0(\mul_a1/fa1_c2_r[14] ), 
        .CI(\mul_a1/fa1_s2_r[15] ), .CO(n371), .S0(n362) );
  HS65_GSS_XOR2X3 U338 ( .A(\mul_a1/fa1_s0_r[15] ), .B(\mul_a1/fa1_s1_r[15] ), 
        .Z(n361) );
  HS65_GS_AND2X4 U339 ( .A(\mul_a1/fa1_s0_r[14] ), .B(\mul_a1/fa1_s1_r[14] ), 
        .Z(n360) );
  HS65_GS_AND2X4 U340 ( .A(\mul_a1/fa1_s0_r[15] ), .B(\mul_a1/fa1_s1_r[15] ), 
        .Z(n379) );
  HS65_GSS_XOR2X3 U341 ( .A(\mul_a1/fa1_s0_r[16] ), .B(\mul_a1/fa1_s1_r[16] ), 
        .Z(n377) );
  HS65_GSS_XOR2X3 U342 ( .A(\mul_a1/fa1_s0_r[12] ), .B(\mul_a1/fa1_s1_r[12] ), 
        .Z(n320) );
  HS65_GS_AND2X4 U343 ( .A(\mul_a1/fa1_s0_r[11] ), .B(\mul_a1/fa1_s1_r[11] ), 
        .Z(n319) );
  HS65_GS_AND2X4 U344 ( .A(\mul_a1/fa1_s0_r[12] ), .B(\mul_a1/fa1_s1_r[12] ), 
        .Z(n356) );
  HS65_GSS_XOR2X3 U345 ( .A(\mul_a1/fa1_c1_r[12] ), .B(\mul_a1/fa1_s2_r[13] ), 
        .Z(n355) );
  HS65_GSS_XOR2X3 U346 ( .A(\mul_a1/fa1_s0_r[13] ), .B(\mul_a1/fa1_s1_r[13] ), 
        .Z(n354) );
  HS65_GS_AND2X4 U347 ( .A(n349), .B(n350), .Z(n598) );
  HS65_GS_FA1X4 U348 ( .A0(\mul_a1/fa1_c1_r[11] ), .B0(n320), .CI(n319), .CO(
        n349), .S0(n347) );
  HS65_GSS_XOR2X3 U349 ( .A(\mul_a1/fa1_s0_r[11] ), .B(\mul_a1/fa1_s1_r[11] ), 
        .Z(n322) );
  HS65_GS_AND2X4 U350 ( .A(\mul_a1/fa1_s0_r[10] ), .B(\mul_a1/fa1_s1_r[10] ), 
        .Z(n321) );
  HS65_GSS_XOR2X3 U351 ( .A(n347), .B(n348), .Z(n346) );
  HS65_GSS_XOR2X3 U352 ( .A(\mul_a1/fa1_s0_r[10] ), .B(\mul_a1/fa1_s1_r[10] ), 
        .Z(n324) );
  HS65_GS_AND2X4 U353 ( .A(\mul_a1/fa1_s0_r[9] ), .B(\mul_a1/fa1_s1_r[9] ), 
        .Z(n323) );
  HS65_GS_FA1X4 U354 ( .A0(\mul_a1/fa1_c1_r[10] ), .B0(n322), .CI(n321), .CO(
        n348), .S0(n327) );
  HS65_GS_AND2X4 U355 ( .A(n326), .B(n327), .Z(n345) );
  HS65_GSS_XOR2X3 U356 ( .A(\mul_a1/fa1_s0_r[9] ), .B(\mul_a1/fa1_s1_r[9] ), 
        .Z(n330) );
  HS65_GS_AND2X4 U357 ( .A(\mul_a1/fa1_s0_r[8] ), .B(\mul_a1/fa1_s1_r[8] ), 
        .Z(n329) );
  HS65_GS_FA1X4 U358 ( .A0(\mul_a1/fa1_c1_r[9] ), .B0(n324), .CI(n323), .CO(
        n326), .S0(n340) );
  HS65_GS_AND2X4 U359 ( .A(n325), .B(n340), .Z(n343) );
  HS65_GSS_XOR2X3 U360 ( .A(n327), .B(n326), .Z(n342) );
  HS65_GSS_XOR2X3 U361 ( .A(\mul_a1/fa1_s0_r[8] ), .B(\mul_a1/fa1_s1_r[8] ), 
        .Z(n334) );
  HS65_GS_AND2X4 U362 ( .A(\mul_a1/fa1_s0_r[7] ), .B(\mul_a1/fa1_s1_r[7] ), 
        .Z(n328) );
  HS65_GS_AND2X4 U363 ( .A(n334), .B(n328), .Z(n331) );
  HS65_GS_FA1X4 U364 ( .A0(\mul_a1/fa1_c1_r[8] ), .B0(n330), .CI(n329), .CO(
        n325), .S0(n336) );
  HS65_GS_AND2X4 U365 ( .A(n331), .B(n336), .Z(n339) );
  HS65_GS_AND2X4 U366 ( .A(\mul_a1/fa1_s0_r[6] ), .B(\mul_a1/fa1_s1_r[6] ), 
        .Z(n333) );
  HS65_GSS_XOR2X3 U367 ( .A(\mul_a1/fa1_s0_r[7] ), .B(\mul_a1/fa1_s1_r[7] ), 
        .Z(n332) );
  HS65_GS_AND2X4 U368 ( .A(n333), .B(n332), .Z(n335) );
  HS65_GS_AND2X4 U369 ( .A(n335), .B(n334), .Z(n337) );
  HS65_GS_AND2X4 U370 ( .A(n337), .B(n336), .Z(n338) );
  HS65_GS_PAO2X4 U371 ( .A(n340), .B(n339), .P(n338), .Z(n341) );
  HS65_GS_PAO2X4 U372 ( .A(n343), .B(n342), .P(n341), .Z(n344) );
  HS65_GS_PAO2X4 U373 ( .A(n346), .B(n345), .P(n344), .Z(n353) );
  HS65_GS_AND2X4 U374 ( .A(n348), .B(n347), .Z(n352) );
  HS65_GSS_XOR2X3 U375 ( .A(n350), .B(n349), .Z(n351) );
  HS65_GS_PAO2X4 U376 ( .A(n353), .B(n352), .P(n351), .Z(n597) );
  HS65_GS_FA1X4 U377 ( .A0(n356), .B0(n355), .CI(n354), .CO(n365), .S0(n350)
         );
  HS65_GS_AND2X4 U378 ( .A(\mul_a1/fa1_c1_r[12] ), .B(\mul_a1/fa1_s2_r[13] ), 
        .Z(n364) );
  HS65_GS_AND2X4 U379 ( .A(\mul_a1/fa1_s0_r[13] ), .B(\mul_a1/fa1_s1_r[13] ), 
        .Z(n359) );
  HS65_GSS_XOR2X3 U380 ( .A(\mul_a1/fa1_s2_r[14] ), .B(\mul_a1/fa1_c1_r[13] ), 
        .Z(n358) );
  HS65_GSS_XOR2X3 U381 ( .A(\mul_a1/fa1_s0_r[14] ), .B(\mul_a1/fa1_s1_r[14] ), 
        .Z(n357) );
  HS65_GS_AND2X4 U382 ( .A(\mul_a1/fa1_c1_r[13] ), .B(\mul_a1/fa1_s2_r[14] ), 
        .Z(n368) );
  HS65_GS_FA1X4 U383 ( .A0(n359), .B0(n358), .CI(n357), .CO(n367), .S0(n363)
         );
  HS65_GS_FA1X4 U384 ( .A0(n362), .B0(n361), .CI(n360), .CO(n370), .S0(n366)
         );
  HS65_GS_FA1X4 U385 ( .A0(n365), .B0(n364), .CI(n363), .CO(n619), .S0(n596)
         );
  HS65_GS_FA1X4 U386 ( .A0(n368), .B0(n367), .CI(n366), .CO(n624), .S0(n620)
         );
  HS65_GS_FA1X4 U387 ( .A0(n371), .B0(n370), .CI(n369), .CO(n373), .S0(n623)
         );
  HS65_GS_NOR2X2 U388 ( .A(n372), .B(n373), .Z(n380) );
  HS65_GS_AOI12X2 U389 ( .A(n373), .B(n372), .C(n380), .Z(n627) );
  HS65_GS_FA1X4 U390 ( .A0(n376), .B0(n375), .CI(n374), .CO(n386), .S0(n384)
         );
  HS65_GS_FA1X4 U391 ( .A0(\mul_a1/fa1_c1_r[15] ), .B0(\mul_a1/fa1_c2_r[15] ), 
        .CI(\mul_a1/fa1_s2_r[16] ), .CO(n383), .S0(n378) );
  HS65_GS_FA1X4 U392 ( .A0(n379), .B0(n378), .CI(n377), .CO(n382), .S0(n369)
         );
  HS65_GS_IVX2 U393 ( .A(n628), .Z(n381) );
  HS65_GS_AOI12X2 U394 ( .A(n627), .B(n381), .C(n380), .Z(n632) );
  HS65_GS_FA1X4 U395 ( .A0(n384), .B0(n383), .CI(n382), .CO(n631), .S0(n628)
         );
  HS65_GS_FA1X4 U396 ( .A0(n387), .B0(n386), .CI(n385), .CO(n636), .S0(n630)
         );
  HS65_GS_FA1X4 U397 ( .A0(n390), .B0(n389), .CI(n388), .CO(n640), .S0(n634)
         );
  HS65_GS_FA1X4 U398 ( .A0(n393), .B0(n392), .CI(n391), .CO(n644), .S0(n638)
         );
  HS65_GS_FA1X4 U399 ( .A0(n396), .B0(n395), .CI(n394), .CO(n648), .S0(n642)
         );
  HS65_GS_FA1X4 U400 ( .A0(n399), .B0(n398), .CI(n397), .CO(n652), .S0(n646)
         );
  HS65_GS_FA1X4 U401 ( .A0(n402), .B0(n401), .CI(n400), .CO(n656), .S0(n650)
         );
  HS65_GS_FA1X4 U402 ( .A0(n405), .B0(n404), .CI(n403), .CO(n660), .S0(n654)
         );
  HS65_GS_FA1X4 U403 ( .A0(n408), .B0(n407), .CI(n406), .CO(n664), .S0(n658)
         );
  HS65_GS_FA1X4 U404 ( .A0(n411), .B0(n410), .CI(n409), .CO(n668), .S0(n662)
         );
  HS65_GS_FA1X4 U405 ( .A0(n414), .B0(n413), .CI(n412), .CO(n672), .S0(n666)
         );
  HS65_GS_FA1X4 U406 ( .A0(n417), .B0(n416), .CI(n415), .CO(n605), .S0(n670)
         );
  HS65_GS_FA1X4 U407 ( .A0(n420), .B0(n419), .CI(n418), .CO(n601), .S0(n603)
         );
  HS65_GS_AND2X4 U408 ( .A(\mul_a1/fa1_s0_r[29] ), .B(\mul_a1/fa1_s1_r[29] ), 
        .Z(n429) );
  HS65_GSS_XOR2X3 U409 ( .A(\mul_a1/fa1_s0_r[30] ), .B(\mul_a1/fa1_s1_r[30] ), 
        .Z(n427) );
  HS65_GS_FA1X4 U410 ( .A0(\mul_a1/fa1_c1_r[28] ), .B0(\mul_a1/fa1_c2_r[28] ), 
        .CI(\mul_a1/fa1_s2_r[29] ), .CO(n425), .S0(n422) );
  HS65_GS_FA1X4 U411 ( .A0(n423), .B0(n422), .CI(n421), .CO(n424), .S0(n418)
         );
  HS65_GS_FA1X4 U412 ( .A0(n426), .B0(n425), .CI(n424), .CO(n607), .S0(n599)
         );
  HS65_GS_FA1X4 U413 ( .A0(\mul_a1/fa1_c1_r[29] ), .B0(\mul_a1/fa1_c2_r[29] ), 
        .CI(\mul_a1/fa1_s2_r[30] ), .CO(n435), .S0(n428) );
  HS65_GS_FA1X4 U414 ( .A0(n429), .B0(n428), .CI(n427), .CO(n434), .S0(n426)
         );
  HS65_GS_AND2X4 U415 ( .A(\mul_a1/fa1_s0_r[30] ), .B(\mul_a1/fa1_s1_r[30] ), 
        .Z(n432) );
  HS65_GSS_XOR2X3 U416 ( .A(\mul_a1/fa1_s2_r[31] ), .B(\mul_a1/fa1_c1_r[30] ), 
        .Z(n431) );
  HS65_GSS_XOR2X3 U417 ( .A(\mul_a1/fa1_s0_r[31] ), .B(\mul_a1/fa1_s1_r[31] ), 
        .Z(n430) );
  HS65_GS_AND2X4 U418 ( .A(\mul_a1/fa1_c1_r[30] ), .B(\mul_a1/fa1_s2_r[31] ), 
        .Z(n438) );
  HS65_GS_FA1X4 U419 ( .A0(n432), .B0(n431), .CI(n430), .CO(n437), .S0(n433)
         );
  HS65_GS_AND2X4 U420 ( .A(\mul_a1/fa1_s0_r[31] ), .B(\mul_a1/fa1_s1_r[31] ), 
        .Z(n441) );
  HS65_GS_NAND2X2 U421 ( .A(\mul_a1/fa1_s0_r[32] ), .B(\mul_a1/fa1_s1_r[32] ), 
        .Z(n444) );
  HS65_GS_OA12X4 U422 ( .A(\mul_a1/fa1_s0_r[32] ), .B(\mul_a1/fa1_s1_r[32] ), 
        .C(n444), .Z(n440) );
  HS65_GSS_XOR2X3 U423 ( .A(\mul_a1/fa1_s2_r[32] ), .B(\mul_a1/fa1_c1_r[31] ), 
        .Z(n439) );
  HS65_GS_FA1X4 U424 ( .A0(n435), .B0(n434), .CI(n433), .CO(n609), .S0(n606)
         );
  HS65_GS_FA1X4 U425 ( .A0(n438), .B0(n437), .CI(n436), .CO(n443), .S0(n610)
         );
  HS65_GS_FA1X4 U426 ( .A0(n441), .B0(n440), .CI(n439), .CO(n442), .S0(n436)
         );
  HS65_GSS_XOR3X2 U427 ( .A(n443), .B(\mul_a1/fa1_s1_r[33] ), .C(n442), .Z(
        n446) );
  HS65_GS_IVX2 U428 ( .A(n444), .Z(n445) );
  HS65_GSS_XOR3X2 U429 ( .A(n447), .B(n446), .C(n445), .Z(n448) );
  HS65_GSS_XOR3X2 U430 ( .A(\mul_a1/fa1_s0_r[33] ), .B(\mul_a1/fa1_c1_r[32] ), 
        .C(n448), .Z(n449) );
  HS65_GSS_XOR3X2 U431 ( .A(n450), .B(\mul_a1/fa1_s2_r[33] ), .C(n449), .Z(
        \mul_a1/result_sat[15] ) );
  HS65_GSS_XOR2X3 U432 ( .A(y_z1[1]), .B(\mul_a1/fa1_s2[13] ), .Z(
        \mul_a1/fa1_s2[14] ) );
  HS65_GS_IVX2 U433 ( .A(y_z1[15]), .Z(n767) );
  HS65_GS_IVX2 U434 ( .A(n767), .Z(\DP_OP_426J1_214_8117/n94 ) );
  HS65_GS_IVX2 U435 ( .A(x_z2[15]), .Z(n1030) );
  HS65_GS_IVX2 U436 ( .A(x_z2[14]), .Z(n1029) );
  HS65_GS_IVX2 U437 ( .A(x_z2[13]), .Z(n1028) );
  HS65_GS_IVX2 U438 ( .A(x_z2[12]), .Z(n1027) );
  HS65_GS_IVX2 U439 ( .A(x_z2[11]), .Z(n1026) );
  HS65_GS_IVX2 U440 ( .A(x_z2[10]), .Z(n1025) );
  HS65_GS_IVX2 U441 ( .A(x_z2[9]), .Z(n1024) );
  HS65_GS_IVX2 U442 ( .A(x_z2[7]), .Z(n1023) );
  HS65_GS_IVX2 U443 ( .A(x_z2[6]), .Z(n1022) );
  HS65_GS_IVX2 U444 ( .A(x_z2[5]), .Z(n1021) );
  HS65_GS_IVX2 U445 ( .A(x_z2[4]), .Z(n1020) );
  HS65_GS_IVX2 U446 ( .A(x_z2[3]), .Z(n1019) );
  HS65_GS_IVX2 U447 ( .A(x_z2[2]), .Z(n1018) );
  HS65_GS_IVX2 U448 ( .A(x_z2[1]), .Z(n1017) );
  HS65_GS_IVX2 U449 ( .A(\mul_b1/fa1_s1[7] ), .Z(n1016) );
  HS65_GS_HA1X4 U450 ( .A0(n1017), .B0(n1016), .CO(n451) );
  HS65_GS_HA1X4 U451 ( .A0(n1018), .B0(n451), .CO(n1012) );
  HS65_GS_NOR2X5 U452 ( .A(x_z2[15]), .B(n957), .Z(n1051) );
  HS65_GS_IVX2 U453 ( .A(y_z1[1]), .Z(n1015) );
  HS65_GS_IVX2 U454 ( .A(\mul_a1/fa1_s2[13] ), .Z(n1014) );
  HS65_GSS_XOR2X3 U455 ( .A(y_z1[2]), .B(n751), .Z(\mul_a1/fa1_s2[15] ) );
  HS65_GS_IVX2 U456 ( .A(y_z1[2]), .Z(n685) );
  HS65_GS_HA1X4 U457 ( .A0(n1015), .B0(n1014), .CO(n452), .S0(n751) );
  HS65_GSS_XOR2X3 U458 ( .A(y_z1[3]), .B(n752), .Z(\mul_a1/fa1_s2[16] ) );
  HS65_GS_IVX2 U459 ( .A(y_z1[3]), .Z(n688) );
  HS65_GS_HA1X4 U460 ( .A0(n685), .B0(n452), .CO(n453), .S0(n752) );
  HS65_GSS_XOR2X3 U461 ( .A(y_z1[4]), .B(n753), .Z(\mul_a1/fa1_s2[17] ) );
  HS65_GS_IVX2 U462 ( .A(y_z1[4]), .Z(n691) );
  HS65_GS_HA1X4 U463 ( .A0(n688), .B0(n453), .CO(n454), .S0(n753) );
  HS65_GSS_XOR2X3 U464 ( .A(y_z1[5]), .B(n754), .Z(\mul_a1/fa1_s2[18] ) );
  HS65_GS_IVX2 U465 ( .A(y_z1[5]), .Z(n694) );
  HS65_GS_HA1X4 U466 ( .A0(n691), .B0(n454), .CO(n455), .S0(n754) );
  HS65_GSS_XOR2X3 U467 ( .A(y_z1[6]), .B(n755), .Z(\mul_a1/fa1_s2[19] ) );
  HS65_GS_IVX2 U468 ( .A(y_z1[6]), .Z(n698) );
  HS65_GS_HA1X4 U469 ( .A0(n694), .B0(n455), .CO(n456), .S0(n755) );
  HS65_GSS_XOR2X3 U470 ( .A(y_z1[7]), .B(n756), .Z(\mul_a1/fa1_s2[20] ) );
  HS65_GS_IVX2 U471 ( .A(y_z1[7]), .Z(n701) );
  HS65_GS_HA1X4 U472 ( .A0(n698), .B0(n456), .CO(n457), .S0(n756) );
  HS65_GSS_XOR2X3 U473 ( .A(y_z1[8]), .B(n757), .Z(\mul_a1/fa1_s2[21] ) );
  HS65_GS_IVX2 U474 ( .A(y_z1[8]), .Z(n704) );
  HS65_GS_HA1X4 U475 ( .A0(n701), .B0(n457), .CO(n458), .S0(n757) );
  HS65_GSS_XOR2X3 U476 ( .A(y_z1[9]), .B(n758), .Z(\mul_a1/fa1_s2[22] ) );
  HS65_GS_IVX2 U477 ( .A(y_z1[9]), .Z(n708) );
  HS65_GS_HA1X4 U478 ( .A0(n704), .B0(n458), .CO(n459), .S0(n758) );
  HS65_GSS_XOR2X3 U479 ( .A(y_z1[10]), .B(n759), .Z(\mul_a1/fa1_s2[23] ) );
  HS65_GS_IVX2 U480 ( .A(y_z1[10]), .Z(n712) );
  HS65_GS_HA1X4 U481 ( .A0(n708), .B0(n459), .CO(n460), .S0(n759) );
  HS65_GSS_XOR2X3 U482 ( .A(y_z1[11]), .B(n760), .Z(\mul_a1/fa1_s2[24] ) );
  HS65_GS_IVX2 U483 ( .A(y_z1[11]), .Z(n715) );
  HS65_GS_HA1X4 U484 ( .A0(n712), .B0(n460), .CO(n461), .S0(n760) );
  HS65_GSS_XOR2X3 U485 ( .A(y_z1[12]), .B(n761), .Z(\mul_a1/fa1_s2[25] ) );
  HS65_GS_IVX2 U486 ( .A(y_z1[12]), .Z(n718) );
  HS65_GS_HA1X4 U487 ( .A0(n715), .B0(n461), .CO(n462), .S0(n761) );
  HS65_GSS_XOR2X3 U488 ( .A(y_z1[13]), .B(n762), .Z(\mul_a1/fa1_s2[26] ) );
  HS65_GS_IVX2 U489 ( .A(y_z1[13]), .Z(n706) );
  HS65_GS_HA1X4 U490 ( .A0(n718), .B0(n462), .CO(n676), .S0(n762) );
  HS65_GSS_XOR2X3 U491 ( .A(y_z1[14]), .B(n763), .Z(\mul_a1/fa1_s2[27] ) );
  HS65_GS_IVX2 U492 ( .A(n463), .Z(n744) );
  HS65_GS_IVX2 U493 ( .A(y_z1[14]), .Z(n710) );
  HS65_GS_HA1X4 U494 ( .A0(n706), .B0(n464), .CO(n466), .S0(n463) );
  HS65_GS_IVX2 U495 ( .A(n465), .Z(n745) );
  HS65_GS_HA1X4 U496 ( .A0(n710), .B0(n466), .CO(n468), .S0(n465) );
  HS65_GS_OR2X4 U497 ( .A(\DP_OP_426J1_214_8117/n94 ), .B(n747), .Z(n749) );
  HS65_GS_IVX2 U498 ( .A(n749), .Z(\mul_a1/fa1_c1[27] ) );
  HS65_GSS_XOR2X3 U499 ( .A(\mul_a1/fa1_s2[13] ), .B(n1010), .Z(
        \mul_a1/fa1_s1[8] ) );
  HS65_GS_HA1X4 U500 ( .A0(n685), .B0(n467), .CO(n469), .S0(n1010) );
  HS65_GSS_XOR2X3 U501 ( .A(y_z1[1]), .B(n1011), .Z(\mul_a1/fa1_s1[9] ) );
  HS65_GS_HA1X4 U502 ( .A0(n767), .B0(n468), .CO(n747), .S0(n1054) );
  HS65_GS_HA1X4 U503 ( .A0(n688), .B0(n469), .CO(n682), .S0(n1011) );
  HS65_GS_NOR2X2 U504 ( .A(\DP_OP_426J1_214_8117/n94 ), .B(n716), .Z(n1052) );
  HS65_GS_IVX2 U505 ( .A(x_z1[15]), .Z(n878) );
  HS65_GS_MUX21I1X3 U506 ( .D0(n878), .D1(data_in[15]), .S0(valid_in), .Z(
        n3464) );
  HS65_GS_IVX2 U507 ( .A(valid_T3), .Z(n1006) );
  HS65_GS_IVX2 U508 ( .A(p_b1[15]), .Z(n502) );
  HS65_GS_IVX2 U509 ( .A(p_b0[15]), .Z(n501) );
  HS65_GS_NAND2X2 U510 ( .A(p_b0[0]), .B(p_b1[0]), .Z(n488) );
  HS65_GS_IVX2 U511 ( .A(n488), .Z(n489) );
  HS65_GS_NAND2X2 U512 ( .A(n504), .B(p_a1[15]), .Z(n499) );
  HS65_GS_NOR3X1 U513 ( .A(p_b1[15]), .B(p_b0[15]), .C(n499), .Z(n511) );
  HS65_GS_FA1X4 U514 ( .A0(p_b0[12]), .B0(p_b1[12]), .CI(n470), .CO(n495), 
        .S0(n471) );
  HS65_GS_IVX2 U515 ( .A(n471), .Z(n521) );
  HS65_GS_FA1X4 U516 ( .A0(p_b0[11]), .B0(p_b1[11]), .CI(n472), .CO(n470), 
        .S0(n473) );
  HS65_GS_IVX2 U517 ( .A(n473), .Z(n769) );
  HS65_GS_FA1X4 U518 ( .A0(p_b0[10]), .B0(p_b1[10]), .CI(n474), .CO(n472), 
        .S0(n475) );
  HS65_GS_IVX2 U519 ( .A(n475), .Z(n774) );
  HS65_GS_FA1X4 U520 ( .A0(p_b0[9]), .B0(p_b1[9]), .CI(n476), .CO(n474), .S0(
        n477) );
  HS65_GS_IVX2 U521 ( .A(n477), .Z(n778) );
  HS65_GS_FA1X4 U522 ( .A0(p_b0[8]), .B0(p_b1[8]), .CI(n478), .CO(n476), .S0(
        n479) );
  HS65_GS_IVX2 U523 ( .A(n479), .Z(n525) );
  HS65_GS_FA1X4 U524 ( .A0(p_b0[7]), .B0(p_b1[7]), .CI(n480), .CO(n478), .S0(
        n481) );
  HS65_GS_IVX2 U525 ( .A(n481), .Z(n782) );
  HS65_GS_FA1X4 U526 ( .A0(p_b0[6]), .B0(p_b1[6]), .CI(n482), .CO(n480), .S0(
        n483) );
  HS65_GS_IVX2 U527 ( .A(n483), .Z(n786) );
  HS65_GS_FA1X4 U528 ( .A0(p_b0[5]), .B0(p_b1[5]), .CI(n484), .CO(n482), .S0(
        n485) );
  HS65_GS_IVX2 U529 ( .A(n485), .Z(n1004) );
  HS65_GS_FA1X4 U530 ( .A0(p_b0[4]), .B0(p_b1[4]), .CI(n486), .CO(n484), .S0(
        n487) );
  HS65_GS_IVX2 U531 ( .A(n487), .Z(n997) );
  HS65_GS_OAI21X2 U532 ( .A(p_b0[0]), .B(p_b1[0]), .C(n488), .Z(n1001) );
  HS65_GS_NAND2X2 U533 ( .A(p_a1[0]), .B(n1001), .Z(n1000) );
  HS65_GS_IVX2 U534 ( .A(n1000), .Z(n590) );
  HS65_GS_FA1X4 U535 ( .A0(p_b0[1]), .B0(p_b1[1]), .CI(n489), .CO(n491), .S0(
        n490) );
  HS65_GS_IVX2 U536 ( .A(n490), .Z(n589) );
  HS65_GS_FA1X4 U537 ( .A0(p_b0[2]), .B0(p_b1[2]), .CI(n491), .CO(n493), .S0(
        n492) );
  HS65_GS_IVX2 U538 ( .A(n492), .Z(n585) );
  HS65_GS_FA1X4 U539 ( .A0(p_b0[3]), .B0(p_b1[3]), .CI(n493), .CO(n486), .S0(
        n494) );
  HS65_GS_IVX2 U540 ( .A(n494), .Z(n581) );
  HS65_GS_FA1X4 U541 ( .A0(p_b0[13]), .B0(p_b1[13]), .CI(n495), .CO(n497), 
        .S0(n496) );
  HS65_GS_IVX2 U542 ( .A(n496), .Z(n516) );
  HS65_GS_FA1X4 U543 ( .A0(p_b0[14]), .B0(p_b1[14]), .CI(n497), .CO(n500), 
        .S0(n498) );
  HS65_GS_IVX2 U544 ( .A(n498), .Z(n506) );
  HS65_GS_OAI21X2 U545 ( .A(n504), .B(p_a1[15]), .C(n499), .Z(n508) );
  HS65_GS_FA1X4 U546 ( .A0(n502), .B0(n501), .CI(n500), .CO(n503), .S0(n504)
         );
  HS65_GS_AOI12X2 U547 ( .A(p_a1[15]), .B(n504), .C(n503), .Z(n510) );
  HS65_GS_AOI12X2 U548 ( .A(n509), .B(n508), .C(n510), .Z(n505) );
  HS65_GS_IVX2 U549 ( .A(data_out[15]), .Z(n766) );
  HS65_GS_OAI32X2 U550 ( .A(n1006), .B(n511), .C(n505), .D(valid_T3), .E(n766), 
        .Z(n3416) );
  HS65_GS_FA1X4 U551 ( .A0(p_a1[14]), .B0(n507), .CI(n506), .CO(n509), .S0(
        n515) );
  HS65_GS_NOR2X2 U552 ( .A(n509), .B(n508), .Z(n513) );
  HS65_GS_IVX2 U553 ( .A(n510), .Z(n512) );
  HS65_GS_CBI4I1X3 U554 ( .A(n513), .B(n512), .C(n511), .D(valid_T3), .Z(n770)
         );
  HS65_GS_OAI12X3 U555 ( .A(n513), .B(n512), .C(valid_T3), .Z(n1008) );
  HS65_GS_NAND2X2 U556 ( .A(data_out[14]), .B(n1006), .Z(n514) );
  HS65_GS_CBI4I1X3 U557 ( .A(n515), .B(n770), .C(n1008), .D(n514), .Z(n3413)
         );
  HS65_GS_FA1X4 U558 ( .A0(p_a1[13]), .B0(n517), .CI(n516), .CO(n507), .S0(
        n519) );
  HS65_GS_NAND2X2 U559 ( .A(data_out[13]), .B(n1006), .Z(n518) );
  HS65_GS_CBI4I1X3 U560 ( .A(n519), .B(n770), .C(n1008), .D(n518), .Z(n3410)
         );
  HS65_GS_FA1X4 U561 ( .A0(p_a1[12]), .B0(n521), .CI(n520), .CO(n517), .S0(
        n523) );
  HS65_GS_NAND2X2 U562 ( .A(data_out[12]), .B(n1006), .Z(n522) );
  HS65_GS_CBI4I1X3 U563 ( .A(n523), .B(n770), .C(n1008), .D(n522), .Z(n3407)
         );
  HS65_GS_FA1X4 U564 ( .A0(p_a1[8]), .B0(n525), .CI(n524), .CO(n777), .S0(n527) );
  HS65_GS_NAND2X2 U565 ( .A(data_out[8]), .B(n1006), .Z(n526) );
  HS65_GS_CBI4I1X3 U566 ( .A(n527), .B(n770), .C(n1008), .D(n526), .Z(n3395)
         );
  HS65_GSS_XNOR2X3 U567 ( .A(n528), .B(n535), .Z(n542) );
  HS65_GS_FA1X4 U568 ( .A0(n531), .B0(n530), .CI(n529), .CO(n67), .S0(n541) );
  HS65_GS_FA1X4 U569 ( .A0(n534), .B0(n533), .CI(n532), .CO(n529), .S0(n540)
         );
  HS65_GS_AOI12X2 U570 ( .A(n537), .B(n536), .C(n535), .Z(n539) );
  HS65_GS_NAND3X2 U571 ( .A(n541), .B(n540), .C(n539), .Z(n538) );
  HS65_GS_OAI12X3 U572 ( .A(n542), .B(n538), .C(\mul_b0/result_sat[15] ), .Z(
        n1045) );
  HS65_GS_OAI21X2 U573 ( .A(n546), .B(n545), .C(n1045), .Z(n544) );
  HS65_GS_NOR3X1 U574 ( .A(n541), .B(n540), .C(n539), .Z(n543) );
  HS65_GS_AOI12X3 U575 ( .A(n543), .B(n542), .C(\mul_b0/result_sat[15] ), .Z(
        n832) );
  HS65_GS_IVX2 U576 ( .A(n832), .Z(n1047) );
  HS65_GS_CBI4I1X3 U577 ( .A(n546), .B(n545), .C(n544), .D(n1047), .Z(
        \mul_b0/result_sat[3] ) );
  HS65_GS_IVX2 U578 ( .A(n878), .Z(n1056) );
  HS65_GSS_XNOR2X3 U579 ( .A(n548), .B(n547), .Z(n570) );
  HS65_GS_FA1X4 U580 ( .A0(n551), .B0(n550), .CI(n549), .CO(n284), .S0(n552)
         );
  HS65_GS_IVX2 U581 ( .A(n552), .Z(n567) );
  HS65_GS_FA1X4 U582 ( .A0(n555), .B0(n554), .CI(n553), .CO(n551), .S0(n565)
         );
  HS65_GS_FA1X4 U583 ( .A0(n558), .B0(n557), .CI(n556), .CO(n560), .S0(n564)
         );
  HS65_GS_FA1X4 U584 ( .A0(n561), .B0(n560), .CI(n559), .CO(n554), .S0(n563)
         );
  HS65_GS_NAND3X2 U585 ( .A(n565), .B(n564), .C(n563), .Z(n562) );
  HS65_GS_OAI12X3 U586 ( .A(n567), .B(n562), .C(\mul_b1/result_sat[15] ), .Z(
        n1036) );
  HS65_GS_OAI21X2 U587 ( .A(n569), .B(n570), .C(n1036), .Z(n568) );
  HS65_GS_NOR3X1 U588 ( .A(n565), .B(n564), .C(n563), .Z(n566) );
  HS65_GS_AOI12X3 U589 ( .A(n567), .B(n566), .C(\mul_b1/result_sat[15] ), .Z(
        n933) );
  HS65_GS_IVX2 U590 ( .A(n933), .Z(n1039) );
  HS65_GS_CBI4I1X3 U591 ( .A(n570), .B(n569), .C(n568), .D(n1039), .Z(
        \mul_b1/result_sat[5] ) );
  HS65_GS_NAND2X2 U592 ( .A(n573), .B(n572), .Z(n571) );
  HS65_GS_OAI21X2 U593 ( .A(n573), .B(n572), .C(n571), .Z(n577) );
  HS65_GS_IVX2 U594 ( .A(n574), .Z(n576) );
  HS65_GS_OAI21X2 U595 ( .A(n576), .B(n577), .C(n1045), .Z(n575) );
  HS65_GS_CBI4I1X3 U596 ( .A(n577), .B(n576), .C(n575), .D(n1047), .Z(
        \mul_b0/result_sat[2] ) );
  HS65_GS_IVX2 U597 ( .A(n1030), .Z(n1055) );
  HS65_GS_NOR2X2 U598 ( .A(n1016), .B(n1017), .Z(\mul_b1/fa1_c1[8] ) );
  HS65_GS_NOR2X2 U599 ( .A(n1017), .B(n1018), .Z(\mul_b1/fa1_c1[9] ) );
  HS65_GS_NOR2X2 U600 ( .A(n1018), .B(n1019), .Z(\mul_b1/fa1_c1[10] ) );
  HS65_GS_NOR2X2 U601 ( .A(n1019), .B(n1020), .Z(\mul_b1/fa1_c1[11] ) );
  HS65_GS_NOR2X2 U602 ( .A(n1020), .B(n1021), .Z(\mul_b1/fa1_c1[12] ) );
  HS65_GS_NOR2X2 U603 ( .A(n1021), .B(n1022), .Z(\mul_b1/fa1_c1[13] ) );
  HS65_GS_NOR2X2 U604 ( .A(n1022), .B(n1023), .Z(\mul_b1/fa1_c1[14] ) );
  HS65_GS_NOR2X2 U605 ( .A(n1023), .B(n950), .Z(\mul_b1/fa1_c1[15] ) );
  HS65_GS_NOR2X2 U606 ( .A(n950), .B(n1024), .Z(\mul_b1/fa1_c1[16] ) );
  HS65_GS_NOR2X2 U607 ( .A(n1024), .B(n1025), .Z(\mul_b1/fa1_c1[17] ) );
  HS65_GS_NOR2X2 U608 ( .A(n1025), .B(n1026), .Z(\mul_b1/fa1_c1[18] ) );
  HS65_GS_NOR2X2 U609 ( .A(n1026), .B(n1027), .Z(\mul_b1/fa1_c1[19] ) );
  HS65_GS_NOR2X2 U610 ( .A(n1027), .B(n1028), .Z(\mul_b1/fa1_c1[20] ) );
  HS65_GS_NOR2X2 U611 ( .A(n1028), .B(n1029), .Z(\mul_b1/fa1_c1[21] ) );
  HS65_GS_NOR2X2 U612 ( .A(n1030), .B(n1029), .Z(\mul_b1/fa1_c1[22] ) );
  HS65_GS_IVX2 U613 ( .A(x_z2[8]), .Z(n950) );
  HS65_GS_IVX2 U614 ( .A(n578), .Z(n989) );
  HS65_GS_HA1X4 U615 ( .A0(n1029), .B0(n579), .CO(n991), .S0(n578) );
  HS65_GS_IVX2 U616 ( .A(n580), .Z(n990) );
  HS65_GS_FA1X4 U617 ( .A0(p_a1[3]), .B0(n582), .CI(n581), .CO(n996), .S0(n584) );
  HS65_GS_NAND2X2 U618 ( .A(data_out[3]), .B(n1006), .Z(n583) );
  HS65_GS_CBI4I1X3 U619 ( .A(n584), .B(n770), .C(n1008), .D(n583), .Z(n3380)
         );
  HS65_GS_FA1X4 U620 ( .A0(p_a1[2]), .B0(n586), .CI(n585), .CO(n582), .S0(n588) );
  HS65_GS_NAND2X2 U621 ( .A(data_out[2]), .B(n1006), .Z(n587) );
  HS65_GS_CBI4I1X3 U622 ( .A(n588), .B(n770), .C(n1008), .D(n587), .Z(n3377)
         );
  HS65_GS_FA1X4 U623 ( .A0(p_a1[1]), .B0(n590), .CI(n589), .CO(n586), .S0(n592) );
  HS65_GS_NAND2X2 U624 ( .A(data_out[1]), .B(n1006), .Z(n591) );
  HS65_GS_CBI4I1X3 U625 ( .A(n592), .B(n770), .C(n1008), .D(n591), .Z(n3374)
         );
  HS65_GS_OAI21X2 U626 ( .A(n595), .B(n594), .C(n1045), .Z(n593) );
  HS65_GS_CBI4I1X3 U627 ( .A(n595), .B(n594), .C(n593), .D(n1047), .Z(
        \mul_b0/result_sat[0] ) );
  HS65_GS_FA1X4 U628 ( .A0(n598), .B0(n597), .CI(n596), .CO(n621), .S0(n618)
         );
  HS65_GS_FA1X4 U629 ( .A0(n601), .B0(n600), .CI(n599), .CO(n608), .S0(n602)
         );
  HS65_GS_IVX2 U630 ( .A(n602), .Z(n616) );
  HS65_GS_FA1X4 U631 ( .A0(n605), .B0(n604), .CI(n603), .CO(n600), .S0(n615)
         );
  HS65_GS_FA1X4 U632 ( .A0(n608), .B0(n607), .CI(n606), .CO(n611), .S0(n614)
         );
  HS65_GS_FA1X4 U633 ( .A0(n611), .B0(n610), .CI(n609), .CO(n447), .S0(n613)
         );
  HS65_GS_NAND3X2 U634 ( .A(n615), .B(n614), .C(n613), .Z(n612) );
  HS65_GS_OAI12X3 U635 ( .A(n616), .B(n612), .C(\mul_a1/result_sat[15] ), .Z(
        n674) );
  HS65_GS_NOR3X1 U636 ( .A(n615), .B(n614), .C(n613), .Z(n617) );
  HS65_GS_AOI12X3 U637 ( .A(n617), .B(n616), .C(\mul_a1/result_sat[15] ), .Z(
        n673) );
  HS65_GS_AO12X4 U638 ( .A(n618), .B(n674), .C(n673), .Z(
        \mul_a1/result_sat[0] ) );
  HS65_GS_FA1X4 U639 ( .A0(n621), .B0(n620), .CI(n619), .CO(n625), .S0(n622)
         );
  HS65_GS_OA12X4 U640 ( .A(n673), .B(n622), .C(n674), .Z(
        \mul_a1/result_sat[1] ) );
  HS65_GS_FA1X4 U641 ( .A0(n625), .B0(n624), .CI(n623), .CO(n372), .S0(n626)
         );
  HS65_GS_OA12X4 U642 ( .A(n673), .B(n626), .C(n674), .Z(
        \mul_a1/result_sat[2] ) );
  HS65_GSS_XOR2X3 U643 ( .A(n628), .B(n627), .Z(n629) );
  HS65_GS_OA12X4 U644 ( .A(n673), .B(n629), .C(n674), .Z(
        \mul_a1/result_sat[3] ) );
  HS65_GS_FA1X4 U645 ( .A0(n632), .B0(n631), .CI(n630), .CO(n635), .S0(n633)
         );
  HS65_GS_AO12X4 U646 ( .A(n633), .B(n674), .C(n673), .Z(
        \mul_a1/result_sat[4] ) );
  HS65_GS_FA1X4 U647 ( .A0(n636), .B0(n635), .CI(n634), .CO(n639), .S0(n637)
         );
  HS65_GS_OA12X4 U648 ( .A(n673), .B(n637), .C(n674), .Z(
        \mul_a1/result_sat[5] ) );
  HS65_GS_FA1X4 U649 ( .A0(n640), .B0(n639), .CI(n638), .CO(n643), .S0(n641)
         );
  HS65_GS_AO12X4 U650 ( .A(n641), .B(n674), .C(n673), .Z(
        \mul_a1/result_sat[6] ) );
  HS65_GS_FA1X4 U651 ( .A0(n644), .B0(n643), .CI(n642), .CO(n647), .S0(n645)
         );
  HS65_GS_OA12X4 U652 ( .A(n673), .B(n645), .C(n674), .Z(
        \mul_a1/result_sat[7] ) );
  HS65_GS_FA1X4 U653 ( .A0(n648), .B0(n647), .CI(n646), .CO(n651), .S0(n649)
         );
  HS65_GS_AO12X4 U654 ( .A(n649), .B(n674), .C(n673), .Z(
        \mul_a1/result_sat[8] ) );
  HS65_GS_FA1X4 U655 ( .A0(n652), .B0(n651), .CI(n650), .CO(n655), .S0(n653)
         );
  HS65_GS_OA12X4 U656 ( .A(n673), .B(n653), .C(n674), .Z(
        \mul_a1/result_sat[9] ) );
  HS65_GS_FA1X4 U657 ( .A0(n656), .B0(n655), .CI(n654), .CO(n659), .S0(n657)
         );
  HS65_GS_AO12X4 U658 ( .A(n657), .B(n674), .C(n673), .Z(
        \mul_a1/result_sat[10] ) );
  HS65_GS_FA1X4 U659 ( .A0(n660), .B0(n659), .CI(n658), .CO(n663), .S0(n661)
         );
  HS65_GS_AO12X4 U660 ( .A(n661), .B(n674), .C(n673), .Z(
        \mul_a1/result_sat[11] ) );
  HS65_GS_FA1X4 U661 ( .A0(n664), .B0(n663), .CI(n662), .CO(n667), .S0(n665)
         );
  HS65_GS_AO12X4 U662 ( .A(n665), .B(n674), .C(n673), .Z(
        \mul_a1/result_sat[12] ) );
  HS65_GS_FA1X4 U663 ( .A0(n668), .B0(n667), .CI(n666), .CO(n671), .S0(n669)
         );
  HS65_GS_AO12X4 U664 ( .A(n669), .B(n674), .C(n673), .Z(
        \mul_a1/result_sat[13] ) );
  HS65_GS_FA1X4 U665 ( .A0(n672), .B0(n671), .CI(n670), .CO(n604), .S0(n675)
         );
  HS65_GS_AO12X4 U666 ( .A(n675), .B(n674), .C(n673), .Z(
        \mul_a1/result_sat[14] ) );
  HS65_GS_HA1X4 U667 ( .A0(n706), .B0(n676), .CO(n677), .S0(n763) );
  HS65_GSS_XNOR2X3 U668 ( .A(n764), .B(n767), .Z(\mul_a1/fa1_s2[28] ) );
  HS65_GS_HA1X4 U669 ( .A0(n710), .B0(n677), .CO(n678), .S0(n764) );
  HS65_GSS_XNOR2X3 U670 ( .A(n765), .B(n767), .Z(\mul_a1/fa1_s2[29] ) );
  HS65_GS_HA1X4 U671 ( .A0(n767), .B0(n678), .CO(n680), .S0(n765) );
  HS65_GSS_XNOR2X3 U672 ( .A(\DP_OP_426J1_214_8117/n94 ), .B(n680), .Z(n679)
         );
  HS65_GSS_XNOR2X3 U673 ( .A(n679), .B(n767), .Z(\mul_a1/fa1_s2[30] ) );
  HS65_GS_NOR2X2 U674 ( .A(\DP_OP_426J1_214_8117/n94 ), .B(n680), .Z(n681) );
  HS65_GSS_XNOR2X3 U675 ( .A(n681), .B(n767), .Z(\mul_a1/fa1_s2[31] ) );
  HS65_GS_HA1X4 U676 ( .A0(n691), .B0(n682), .CO(n683), .S0(n719) );
  HS65_GS_PAO2X4 U677 ( .A(\mul_a1/fa1_s2[13] ), .B(n719), .P(y_z1[2]), .Z(
        \mul_a1/fa1_c1[10] ) );
  HS65_GS_HA1X4 U678 ( .A0(n1015), .B0(n1014), .CO(n684), .S0(n721) );
  HS65_GS_HA1X4 U679 ( .A0(n694), .B0(n683), .CO(n686), .S0(n720) );
  HS65_GS_PAO2X4 U680 ( .A(n721), .B(n720), .P(y_z1[3]), .Z(
        \mul_a1/fa1_c1[11] ) );
  HS65_GS_HA1X4 U681 ( .A0(n685), .B0(n684), .CO(n687), .S0(n723) );
  HS65_GS_HA1X4 U682 ( .A0(n698), .B0(n686), .CO(n689), .S0(n722) );
  HS65_GS_PAO2X4 U683 ( .A(n723), .B(n722), .P(y_z1[4]), .Z(
        \mul_a1/fa1_c1[12] ) );
  HS65_GS_HA1X4 U684 ( .A0(n688), .B0(n687), .CO(n690), .S0(n725) );
  HS65_GS_HA1X4 U685 ( .A0(n701), .B0(n689), .CO(n692), .S0(n724) );
  HS65_GS_PAO2X4 U686 ( .A(n725), .B(n724), .P(y_z1[5]), .Z(
        \mul_a1/fa1_c1[13] ) );
  HS65_GS_HA1X4 U687 ( .A0(n691), .B0(n690), .CO(n693), .S0(n727) );
  HS65_GS_HA1X4 U688 ( .A0(n704), .B0(n692), .CO(n695), .S0(n726) );
  HS65_GS_PAO2X4 U689 ( .A(n727), .B(n726), .P(y_z1[6]), .Z(
        \mul_a1/fa1_c1[14] ) );
  HS65_GS_HA1X4 U690 ( .A0(n694), .B0(n693), .CO(n697), .S0(n729) );
  HS65_GS_HA1X4 U691 ( .A0(n708), .B0(n695), .CO(n696), .S0(n728) );
  HS65_GS_PAO2X4 U692 ( .A(n729), .B(n728), .P(y_z1[7]), .Z(
        \mul_a1/fa1_c1[15] ) );
  HS65_GS_HA1X4 U693 ( .A0(n712), .B0(n696), .CO(n699), .S0(n731) );
  HS65_GS_HA1X4 U694 ( .A0(n698), .B0(n697), .CO(n700), .S0(n730) );
  HS65_GS_PAO2X4 U695 ( .A(n731), .B(n730), .P(y_z1[8]), .Z(
        \mul_a1/fa1_c1[16] ) );
  HS65_GS_HA1X4 U696 ( .A0(n715), .B0(n699), .CO(n702), .S0(n733) );
  HS65_GS_HA1X4 U697 ( .A0(n701), .B0(n700), .CO(n703), .S0(n732) );
  HS65_GS_PAO2X4 U698 ( .A(n733), .B(n732), .P(y_z1[9]), .Z(
        \mul_a1/fa1_c1[17] ) );
  HS65_GS_HA1X4 U699 ( .A0(n718), .B0(n702), .CO(n705), .S0(n735) );
  HS65_GS_HA1X4 U700 ( .A0(n704), .B0(n703), .CO(n707), .S0(n734) );
  HS65_GS_PAO2X4 U701 ( .A(n735), .B(n734), .P(y_z1[10]), .Z(
        \mul_a1/fa1_c1[18] ) );
  HS65_GS_HA1X4 U702 ( .A0(n706), .B0(n705), .CO(n709), .S0(n737) );
  HS65_GS_HA1X4 U703 ( .A0(n708), .B0(n707), .CO(n711), .S0(n736) );
  HS65_GS_PAO2X4 U704 ( .A(n737), .B(n736), .P(y_z1[11]), .Z(
        \mul_a1/fa1_c1[19] ) );
  HS65_GS_HA1X4 U705 ( .A0(n710), .B0(n709), .CO(n713), .S0(n739) );
  HS65_GS_HA1X4 U706 ( .A0(n712), .B0(n711), .CO(n714), .S0(n738) );
  HS65_GS_PAO2X4 U707 ( .A(n739), .B(n738), .P(y_z1[12]), .Z(
        \mul_a1/fa1_c1[20] ) );
  HS65_GS_HA1X4 U708 ( .A0(n767), .B0(n713), .CO(n716), .S0(n741) );
  HS65_GS_HA1X4 U709 ( .A0(n715), .B0(n714), .CO(n717), .S0(n740) );
  HS65_GS_PAO2X4 U710 ( .A(n741), .B(n740), .P(y_z1[13]), .Z(
        \mul_a1/fa1_c1[21] ) );
  HS65_GSS_XNOR2X3 U711 ( .A(\DP_OP_426J1_214_8117/n94 ), .B(n716), .Z(n743)
         );
  HS65_GS_HA1X4 U712 ( .A0(n718), .B0(n717), .CO(n464), .S0(n742) );
  HS65_GS_PAO2X4 U713 ( .A(n743), .B(n742), .P(y_z1[14]), .Z(
        \mul_a1/fa1_c1[22] ) );
  HS65_GSS_XOR3X2 U714 ( .A(y_z1[2]), .B(\mul_a1/fa1_s2[13] ), .C(n719), .Z(
        \mul_a1/fa1_s1[10] ) );
  HS65_GSS_XOR3X2 U715 ( .A(y_z1[3]), .B(n721), .C(n720), .Z(
        \mul_a1/fa1_s1[11] ) );
  HS65_GSS_XOR3X2 U716 ( .A(y_z1[4]), .B(n723), .C(n722), .Z(
        \mul_a1/fa1_s1[12] ) );
  HS65_GSS_XOR3X2 U717 ( .A(y_z1[5]), .B(n725), .C(n724), .Z(
        \mul_a1/fa1_s1[13] ) );
  HS65_GSS_XOR3X2 U718 ( .A(y_z1[6]), .B(n727), .C(n726), .Z(
        \mul_a1/fa1_s1[14] ) );
  HS65_GSS_XOR3X2 U719 ( .A(y_z1[7]), .B(n729), .C(n728), .Z(
        \mul_a1/fa1_s1[15] ) );
  HS65_GSS_XOR3X2 U720 ( .A(y_z1[8]), .B(n731), .C(n730), .Z(
        \mul_a1/fa1_s1[16] ) );
  HS65_GSS_XOR3X2 U721 ( .A(y_z1[9]), .B(n733), .C(n732), .Z(
        \mul_a1/fa1_s1[17] ) );
  HS65_GSS_XOR3X2 U722 ( .A(y_z1[10]), .B(n735), .C(n734), .Z(
        \mul_a1/fa1_s1[18] ) );
  HS65_GSS_XOR3X2 U723 ( .A(y_z1[11]), .B(n737), .C(n736), .Z(
        \mul_a1/fa1_s1[19] ) );
  HS65_GSS_XOR3X2 U724 ( .A(y_z1[12]), .B(n739), .C(n738), .Z(
        \mul_a1/fa1_s1[20] ) );
  HS65_GSS_XOR3X2 U725 ( .A(y_z1[13]), .B(n741), .C(n740), .Z(
        \mul_a1/fa1_s1[21] ) );
  HS65_GSS_XOR3X2 U726 ( .A(n743), .B(y_z1[14]), .C(n742), .Z(
        \mul_a1/fa1_s1[22] ) );
  HS65_GSS_XNOR2X3 U727 ( .A(n1052), .B(n767), .Z(n750) );
  HS65_GSS_XNOR2X3 U728 ( .A(n750), .B(n744), .Z(\mul_a1/fa1_s1[23] ) );
  HS65_GSS_XNOR2X3 U729 ( .A(n750), .B(n745), .Z(\mul_a1/fa1_s1[24] ) );
  HS65_GS_IVX2 U730 ( .A(n1054), .Z(n746) );
  HS65_GSS_XNOR2X3 U731 ( .A(n750), .B(n746), .Z(\mul_a1/fa1_s1[25] ) );
  HS65_GSS_XOR2X3 U732 ( .A(\DP_OP_426J1_214_8117/n94 ), .B(n747), .Z(n748) );
  HS65_GSS_XNOR2X3 U733 ( .A(n750), .B(n748), .Z(\mul_a1/fa1_s1[26] ) );
  HS65_GSS_XNOR2X3 U734 ( .A(n750), .B(n749), .Z(\mul_a1/fa1_s1[28] ) );
  HS65_GS_AND2X4 U735 ( .A(\mul_a1/fa1_s2[13] ), .B(y_z1[1]), .Z(
        \mul_a1/fa1_c2[14] ) );
  HS65_GS_AND2X4 U736 ( .A(n751), .B(y_z1[2]), .Z(\mul_a1/fa1_c2[15] ) );
  HS65_GS_AND2X4 U737 ( .A(n752), .B(y_z1[3]), .Z(\mul_a1/fa1_c2[16] ) );
  HS65_GS_AND2X4 U738 ( .A(n753), .B(y_z1[4]), .Z(\mul_a1/fa1_c2[17] ) );
  HS65_GS_AND2X4 U739 ( .A(n754), .B(y_z1[5]), .Z(\mul_a1/fa1_c2[18] ) );
  HS65_GS_AND2X4 U740 ( .A(n755), .B(y_z1[6]), .Z(\mul_a1/fa1_c2[19] ) );
  HS65_GS_AND2X4 U741 ( .A(n756), .B(y_z1[7]), .Z(\mul_a1/fa1_c2[20] ) );
  HS65_GS_AND2X4 U742 ( .A(n757), .B(y_z1[8]), .Z(\mul_a1/fa1_c2[21] ) );
  HS65_GS_AND2X4 U743 ( .A(n758), .B(y_z1[9]), .Z(\mul_a1/fa1_c2[22] ) );
  HS65_GS_AND2X4 U744 ( .A(n759), .B(y_z1[10]), .Z(\mul_a1/fa1_c2[23] ) );
  HS65_GS_AND2X4 U745 ( .A(n760), .B(y_z1[11]), .Z(\mul_a1/fa1_c2[24] ) );
  HS65_GS_AND2X4 U746 ( .A(n761), .B(y_z1[12]), .Z(\mul_a1/fa1_c2[25] ) );
  HS65_GS_AND2X4 U747 ( .A(n762), .B(y_z1[13]), .Z(\mul_a1/fa1_c2[26] ) );
  HS65_GS_AND2X4 U748 ( .A(y_z1[14]), .B(n763), .Z(\mul_a1/fa1_c2[27] ) );
  HS65_GS_AND2X4 U749 ( .A(\DP_OP_426J1_214_8117/n94 ), .B(n764), .Z(
        \mul_a1/fa1_c2[28] ) );
  HS65_GS_AND2X4 U750 ( .A(\DP_OP_426J1_214_8117/n94 ), .B(n765), .Z(
        \mul_a1/fa1_c2[29] ) );
  HS65_GS_MUX21X4 U751 ( .D0(x_z1[14]), .D1(data_in[14]), .S0(valid_in), .Z(
        n3463) );
  HS65_GS_MUX21X4 U752 ( .D0(x_z1[13]), .D1(data_in[13]), .S0(valid_in), .Z(
        n3462) );
  HS65_GS_MUX21X4 U753 ( .D0(x_z1[12]), .D1(data_in[12]), .S0(valid_in), .Z(
        n3461) );
  HS65_GS_MUX21X4 U754 ( .D0(x_z1[11]), .D1(data_in[11]), .S0(valid_in), .Z(
        n3460) );
  HS65_GS_MUX21X4 U755 ( .D0(x_z1[10]), .D1(data_in[10]), .S0(valid_in), .Z(
        n3459) );
  HS65_GS_MUX21X4 U756 ( .D0(x_z1[9]), .D1(data_in[9]), .S0(valid_in), .Z(
        n3458) );
  HS65_GS_MUX21X4 U757 ( .D0(x_z1[8]), .D1(data_in[8]), .S0(valid_in), .Z(
        n3457) );
  HS65_GS_MUX21X4 U758 ( .D0(x_z1[7]), .D1(data_in[7]), .S0(valid_in), .Z(
        n3456) );
  HS65_GS_MUX21X4 U759 ( .D0(x_z1[6]), .D1(data_in[6]), .S0(valid_in), .Z(
        n3455) );
  HS65_GS_MUX21X4 U760 ( .D0(x_z1[5]), .D1(data_in[5]), .S0(valid_in), .Z(
        n3454) );
  HS65_GS_MUX21X4 U761 ( .D0(x_z1[4]), .D1(data_in[4]), .S0(valid_in), .Z(
        n3453) );
  HS65_GS_MUX21X4 U762 ( .D0(x_z1[3]), .D1(data_in[3]), .S0(valid_in), .Z(
        n3452) );
  HS65_GS_MUX21X4 U763 ( .D0(x_z1[2]), .D1(data_in[2]), .S0(valid_in), .Z(
        n3451) );
  HS65_GS_MUX21X4 U764 ( .D0(x_z1[1]), .D1(data_in[1]), .S0(valid_in), .Z(
        n3450) );
  HS65_GS_MUX21X4 U765 ( .D0(x_z1[0]), .D1(data_in[0]), .S0(valid_in), .Z(
        n3449) );
  HS65_GS_MUXI21X2 U766 ( .D0(n1030), .D1(n878), .S0(valid_in), .Z(n3448) );
  HS65_GS_IVX2 U767 ( .A(x_z1[14]), .Z(n869) );
  HS65_GS_MUXI21X2 U768 ( .D0(n1029), .D1(n869), .S0(valid_in), .Z(n3446) );
  HS65_GS_IVX2 U769 ( .A(x_z1[13]), .Z(n867) );
  HS65_GS_MUXI21X2 U770 ( .D0(n1028), .D1(n867), .S0(valid_in), .Z(n3444) );
  HS65_GS_IVX2 U771 ( .A(x_z1[12]), .Z(n865) );
  HS65_GS_MUXI21X2 U772 ( .D0(n1027), .D1(n865), .S0(valid_in), .Z(n3442) );
  HS65_GS_IVX2 U773 ( .A(x_z1[11]), .Z(n863) );
  HS65_GS_MUXI21X2 U774 ( .D0(n1026), .D1(n863), .S0(valid_in), .Z(n3440) );
  HS65_GS_IVX2 U775 ( .A(x_z1[10]), .Z(n861) );
  HS65_GS_MUXI21X2 U776 ( .D0(n1025), .D1(n861), .S0(valid_in), .Z(n3438) );
  HS65_GS_IVX2 U777 ( .A(x_z1[9]), .Z(n859) );
  HS65_GS_MUXI21X2 U778 ( .D0(n1024), .D1(n859), .S0(valid_in), .Z(n3436) );
  HS65_GS_IVX2 U779 ( .A(x_z1[8]), .Z(n857) );
  HS65_GS_MUXI21X2 U780 ( .D0(n950), .D1(n857), .S0(valid_in), .Z(n3434) );
  HS65_GS_IVX2 U781 ( .A(x_z1[7]), .Z(n855) );
  HS65_GS_MUXI21X2 U782 ( .D0(n1023), .D1(n855), .S0(valid_in), .Z(n3432) );
  HS65_GS_IVX2 U783 ( .A(x_z1[6]), .Z(n853) );
  HS65_GS_MUXI21X2 U784 ( .D0(n1022), .D1(n853), .S0(valid_in), .Z(n3430) );
  HS65_GS_IVX2 U785 ( .A(x_z1[5]), .Z(n843) );
  HS65_GS_MUXI21X2 U786 ( .D0(n1021), .D1(n843), .S0(valid_in), .Z(n3428) );
  HS65_GS_IVX2 U787 ( .A(x_z1[4]), .Z(n841) );
  HS65_GS_MUXI21X2 U788 ( .D0(n1020), .D1(n841), .S0(valid_in), .Z(n3426) );
  HS65_GS_IVX2 U789 ( .A(x_z1[3]), .Z(n839) );
  HS65_GS_MUXI21X2 U790 ( .D0(n1019), .D1(n839), .S0(valid_in), .Z(n3424) );
  HS65_GS_IVX2 U791 ( .A(x_z1[2]), .Z(n837) );
  HS65_GS_MUXI21X2 U792 ( .D0(n1018), .D1(n837), .S0(valid_in), .Z(n3422) );
  HS65_GS_IVX2 U793 ( .A(x_z1[1]), .Z(n835) );
  HS65_GS_MUXI21X2 U794 ( .D0(n1017), .D1(n835), .S0(valid_in), .Z(n3420) );
  HS65_GS_IVX2 U795 ( .A(x_z1[0]), .Z(n834) );
  HS65_GS_MUXI21X2 U796 ( .D0(n1016), .D1(n834), .S0(valid_in), .Z(n3418) );
  HS65_GS_MUXI21X2 U797 ( .D0(n767), .D1(n766), .S0(valid_in), .Z(n3415) );
  HS65_GS_MUX21X4 U798 ( .D0(y_z1[14]), .D1(data_out[14]), .S0(valid_in), .Z(
        n3412) );
  HS65_GS_MUX21X4 U799 ( .D0(y_z1[13]), .D1(data_out[13]), .S0(valid_in), .Z(
        n3409) );
  HS65_GS_MUX21X4 U800 ( .D0(y_z1[12]), .D1(data_out[12]), .S0(valid_in), .Z(
        n3406) );
  HS65_GS_FA1X4 U801 ( .A0(p_a1[11]), .B0(n769), .CI(n768), .CO(n520), .S0(
        n772) );
  HS65_GS_IVX2 U802 ( .A(n770), .Z(n1005) );
  HS65_GS_AOI12X2 U803 ( .A(data_out[11]), .B(n1006), .C(n1005), .Z(n771) );
  HS65_GS_OAI21X2 U804 ( .A(n772), .B(n1008), .C(n771), .Z(n3404) );
  HS65_GS_MUX21X4 U805 ( .D0(y_z1[11]), .D1(data_out[11]), .S0(valid_in), .Z(
        n3403) );
  HS65_GS_FA1X4 U806 ( .A0(p_a1[10]), .B0(n774), .CI(n773), .CO(n768), .S0(
        n776) );
  HS65_GS_AOI12X2 U807 ( .A(data_out[10]), .B(n1006), .C(n1005), .Z(n775) );
  HS65_GS_OAI21X2 U808 ( .A(n776), .B(n1008), .C(n775), .Z(n3401) );
  HS65_GS_MUX21X4 U809 ( .D0(y_z1[10]), .D1(data_out[10]), .S0(valid_in), .Z(
        n3400) );
  HS65_GS_FA1X4 U810 ( .A0(p_a1[9]), .B0(n778), .CI(n777), .CO(n773), .S0(n780) );
  HS65_GS_AOI12X2 U811 ( .A(data_out[9]), .B(n1006), .C(n1005), .Z(n779) );
  HS65_GS_OAI21X2 U812 ( .A(n780), .B(n1008), .C(n779), .Z(n3398) );
  HS65_GS_MUX21X4 U813 ( .D0(y_z1[9]), .D1(data_out[9]), .S0(valid_in), .Z(
        n3397) );
  HS65_GS_MUX21X4 U814 ( .D0(y_z1[8]), .D1(data_out[8]), .S0(valid_in), .Z(
        n3394) );
  HS65_GS_FA1X4 U815 ( .A0(p_a1[7]), .B0(n782), .CI(n781), .CO(n524), .S0(n784) );
  HS65_GS_AOI12X2 U816 ( .A(data_out[7]), .B(n1006), .C(n1005), .Z(n783) );
  HS65_GS_OAI21X2 U817 ( .A(n784), .B(n1008), .C(n783), .Z(n3392) );
  HS65_GS_MUX21X4 U818 ( .D0(y_z1[7]), .D1(data_out[7]), .S0(valid_in), .Z(
        n3391) );
  HS65_GS_FA1X4 U819 ( .A0(p_a1[6]), .B0(n786), .CI(n785), .CO(n781), .S0(n788) );
  HS65_GS_AOI12X2 U820 ( .A(data_out[6]), .B(n1006), .C(n1005), .Z(n787) );
  HS65_GS_OAI21X2 U821 ( .A(n788), .B(n1008), .C(n787), .Z(n3389) );
  HS65_GS_MUX21X4 U822 ( .D0(y_z1[6]), .D1(data_out[6]), .S0(valid_in), .Z(
        n3388) );
  HS65_GS_FA1X4 U823 ( .A0(n791), .B0(n790), .CI(n789), .CO(n793), .S0(n792)
         );
  HS65_GS_OA12X4 U824 ( .A(n832), .B(n792), .C(n1045), .Z(
        \mul_b0/result_sat[4] ) );
  HS65_GS_FA1X4 U825 ( .A0(n795), .B0(n794), .CI(n793), .CO(n797), .S0(n796)
         );
  HS65_GS_AO12X4 U826 ( .A(n796), .B(n1045), .C(n832), .Z(
        \mul_b0/result_sat[5] ) );
  HS65_GS_FA1X4 U827 ( .A0(n799), .B0(n798), .CI(n797), .CO(n801), .S0(n800)
         );
  HS65_GS_OA12X4 U828 ( .A(n832), .B(n800), .C(n1045), .Z(
        \mul_b0/result_sat[6] ) );
  HS65_GS_FA1X4 U829 ( .A0(n803), .B0(n802), .CI(n801), .CO(n807), .S0(n804)
         );
  HS65_GS_AO12X4 U830 ( .A(n804), .B(n1045), .C(n832), .Z(
        \mul_b0/result_sat[7] ) );
  HS65_GS_FA1X4 U831 ( .A0(n807), .B0(n806), .CI(n805), .CO(n811), .S0(n808)
         );
  HS65_GS_AO12X4 U832 ( .A(n808), .B(n1045), .C(n832), .Z(
        \mul_b0/result_sat[8] ) );
  HS65_GS_FA1X4 U833 ( .A0(n811), .B0(n810), .CI(n809), .CO(n813), .S0(n812)
         );
  HS65_GS_AO12X4 U834 ( .A(n812), .B(n1045), .C(n832), .Z(
        \mul_b0/result_sat[9] ) );
  HS65_GS_FA1X4 U835 ( .A0(n815), .B0(n814), .CI(n813), .CO(n817), .S0(n816)
         );
  HS65_GS_OA12X4 U836 ( .A(n832), .B(n816), .C(n1045), .Z(
        \mul_b0/result_sat[10] ) );
  HS65_GS_FA1X4 U837 ( .A0(n819), .B0(n818), .CI(n817), .CO(n823), .S0(n820)
         );
  HS65_GS_AO12X4 U838 ( .A(n820), .B(n1045), .C(n832), .Z(
        \mul_b0/result_sat[11] ) );
  HS65_GS_FA1X4 U839 ( .A0(n823), .B0(n822), .CI(n821), .CO(n827), .S0(n824)
         );
  HS65_GS_AO12X4 U840 ( .A(n824), .B(n1045), .C(n832), .Z(
        \mul_b0/result_sat[12] ) );
  HS65_GS_FA1X4 U841 ( .A0(n827), .B0(n826), .CI(n825), .CO(n831), .S0(n828)
         );
  HS65_GS_AO12X4 U842 ( .A(n828), .B(n1045), .C(n832), .Z(
        \mul_b0/result_sat[13] ) );
  HS65_GS_FA1X4 U843 ( .A0(n831), .B0(n830), .CI(n829), .CO(n532), .S0(n833)
         );
  HS65_GS_AO12X4 U844 ( .A(n833), .B(n1045), .C(n832), .Z(
        \mul_b0/result_sat[14] ) );
  HS65_GS_AND2X4 U845 ( .A(x_z1[5]), .B(x_z1[0]), .Z(\mul_b0/fa1_c0[5] ) );
  HS65_GS_AND2X4 U846 ( .A(x_z1[6]), .B(n854), .Z(\mul_b0/fa1_c0[6] ) );
  HS65_GS_HA1X4 U847 ( .A0(n835), .B0(n834), .CO(n836), .S0(n854) );
  HS65_GS_AND2X4 U848 ( .A(n856), .B(x_z1[7]), .Z(\mul_b0/fa1_c0[7] ) );
  HS65_GS_HA1X4 U849 ( .A0(n837), .B0(n836), .CO(n838), .S0(n856) );
  HS65_GS_AND2X4 U850 ( .A(x_z1[8]), .B(n858), .Z(\mul_b0/fa1_c0[8] ) );
  HS65_GS_HA1X4 U851 ( .A0(n839), .B0(n838), .CO(n840), .S0(n858) );
  HS65_GS_AND2X4 U852 ( .A(n860), .B(x_z1[9]), .Z(\mul_b0/fa1_c0[9] ) );
  HS65_GS_HA1X4 U853 ( .A0(n841), .B0(n840), .CO(n842), .S0(n860) );
  HS65_GS_AND2X4 U854 ( .A(n862), .B(x_z1[10]), .Z(\mul_b0/fa1_c0[10] ) );
  HS65_GS_HA1X4 U855 ( .A0(n843), .B0(n842), .CO(n844), .S0(n862) );
  HS65_GS_AND2X4 U856 ( .A(n864), .B(x_z1[11]), .Z(\mul_b0/fa1_c0[11] ) );
  HS65_GS_HA1X4 U857 ( .A0(n853), .B0(n844), .CO(n845), .S0(n864) );
  HS65_GS_AND2X4 U858 ( .A(x_z1[12]), .B(n866), .Z(\mul_b0/fa1_c0[12] ) );
  HS65_GS_HA1X4 U859 ( .A0(n855), .B0(n845), .CO(n846), .S0(n866) );
  HS65_GS_AND2X4 U860 ( .A(x_z1[13]), .B(n868), .Z(\mul_b0/fa1_c0[13] ) );
  HS65_GS_HA1X4 U861 ( .A0(n857), .B0(n846), .CO(n847), .S0(n868) );
  HS65_GS_AND2X4 U862 ( .A(x_z1[14]), .B(n870), .Z(\mul_b0/fa1_c0[14] ) );
  HS65_GS_HA1X4 U863 ( .A0(n859), .B0(n847), .CO(n848), .S0(n870) );
  HS65_GS_AND2X4 U864 ( .A(n871), .B(n1056), .Z(\mul_b0/fa1_c0[15] ) );
  HS65_GS_HA1X4 U865 ( .A0(n861), .B0(n848), .CO(n849), .S0(n871) );
  HS65_GS_AND2X4 U866 ( .A(n872), .B(x_z1[15]), .Z(\mul_b0/fa1_c0[16] ) );
  HS65_GS_HA1X4 U867 ( .A0(n863), .B0(n849), .CO(n850), .S0(n872) );
  HS65_GS_AND2X4 U868 ( .A(n873), .B(x_z1[15]), .Z(\mul_b0/fa1_c0[17] ) );
  HS65_GS_HA1X4 U869 ( .A0(n865), .B0(n850), .CO(n851), .S0(n873) );
  HS65_GS_AND2X4 U870 ( .A(n874), .B(x_z1[15]), .Z(\mul_b0/fa1_c0[18] ) );
  HS65_GS_HA1X4 U871 ( .A0(n867), .B0(n851), .CO(n852), .S0(n874) );
  HS65_GS_AND2X4 U872 ( .A(n875), .B(x_z1[15]), .Z(\mul_b0/fa1_c0[19] ) );
  HS65_GS_HA1X4 U873 ( .A0(n869), .B0(n852), .CO(n877), .S0(n875) );
  HS65_GSS_XNOR2X3 U874 ( .A(x_z1[15]), .B(n877), .Z(n876) );
  HS65_GS_AND2X4 U875 ( .A(n876), .B(n1056), .Z(\mul_b0/fa1_c0[20] ) );
  HS65_GSS_XNOR2X3 U876 ( .A(n854), .B(n853), .Z(\mul_b0/fa1_s0[6] ) );
  HS65_GSS_XNOR2X3 U877 ( .A(n856), .B(n855), .Z(\mul_b0/fa1_s0[7] ) );
  HS65_GSS_XNOR2X3 U878 ( .A(n858), .B(n857), .Z(\mul_b0/fa1_s0[8] ) );
  HS65_GSS_XNOR2X3 U879 ( .A(n860), .B(n859), .Z(\mul_b0/fa1_s0[9] ) );
  HS65_GSS_XNOR2X3 U880 ( .A(n862), .B(n861), .Z(\mul_b0/fa1_s0[10] ) );
  HS65_GSS_XNOR2X3 U881 ( .A(n864), .B(n863), .Z(\mul_b0/fa1_s0[11] ) );
  HS65_GSS_XNOR2X3 U882 ( .A(n866), .B(n865), .Z(\mul_b0/fa1_s0[12] ) );
  HS65_GSS_XNOR2X3 U883 ( .A(n868), .B(n867), .Z(\mul_b0/fa1_s0[13] ) );
  HS65_GSS_XNOR2X3 U884 ( .A(n870), .B(n869), .Z(\mul_b0/fa1_s0[14] ) );
  HS65_GSS_XNOR2X3 U885 ( .A(n871), .B(n878), .Z(\mul_b0/fa1_s0[15] ) );
  HS65_GSS_XNOR2X3 U886 ( .A(n872), .B(n878), .Z(\mul_b0/fa1_s0[16] ) );
  HS65_GSS_XNOR2X3 U887 ( .A(n873), .B(n878), .Z(\mul_b0/fa1_s0[17] ) );
  HS65_GSS_XNOR2X3 U888 ( .A(n874), .B(n878), .Z(\mul_b0/fa1_s0[18] ) );
  HS65_GSS_XNOR2X3 U889 ( .A(n875), .B(n878), .Z(\mul_b0/fa1_s0[19] ) );
  HS65_GSS_XNOR2X3 U890 ( .A(n876), .B(n878), .Z(\mul_b0/fa1_s0[20] ) );
  HS65_GS_NOR2X2 U891 ( .A(x_z1[15]), .B(n877), .Z(n879) );
  HS65_GSS_XNOR2X3 U892 ( .A(n879), .B(n878), .Z(\mul_b0/fa1_s0[30] ) );
  HS65_GS_FA1X4 U893 ( .A0(n882), .B0(n881), .CI(n880), .CO(n885), .S0(n883)
         );
  HS65_GS_AO12X4 U894 ( .A(n883), .B(n1036), .C(n933), .Z(
        \mul_b1/result_sat[0] ) );
  HS65_GS_FA1X4 U895 ( .A0(n886), .B0(n885), .CI(n884), .CO(n888), .S0(n887)
         );
  HS65_GS_AO12X4 U896 ( .A(n887), .B(n1036), .C(n933), .Z(
        \mul_b1/result_sat[1] ) );
  HS65_GS_FA1X4 U897 ( .A0(n890), .B0(n889), .CI(n888), .CO(n894), .S0(n891)
         );
  HS65_GS_AO12X4 U898 ( .A(n891), .B(n1036), .C(n933), .Z(
        \mul_b1/result_sat[2] ) );
  HS65_GS_FA1X4 U899 ( .A0(n894), .B0(n893), .CI(n892), .CO(n896), .S0(n895)
         );
  HS65_GS_AO12X4 U900 ( .A(n895), .B(n1036), .C(n933), .Z(
        \mul_b1/result_sat[3] ) );
  HS65_GS_FA1X4 U901 ( .A0(n898), .B0(n897), .CI(n896), .CO(n223), .S0(n899)
         );
  HS65_GS_OA12X4 U902 ( .A(n933), .B(n899), .C(n1036), .Z(
        \mul_b1/result_sat[4] ) );
  HS65_GS_FA1X4 U903 ( .A0(n902), .B0(n901), .CI(n900), .CO(n905), .S0(n903)
         );
  HS65_GS_AO12X4 U904 ( .A(n903), .B(n1036), .C(n933), .Z(
        \mul_b1/result_sat[6] ) );
  HS65_GS_FA1X4 U905 ( .A0(n906), .B0(n905), .CI(n904), .CO(n909), .S0(n907)
         );
  HS65_GS_AO12X4 U906 ( .A(n907), .B(n1036), .C(n933), .Z(
        \mul_b1/result_sat[7] ) );
  HS65_GS_FA1X4 U907 ( .A0(n910), .B0(n909), .CI(n908), .CO(n913), .S0(n911)
         );
  HS65_GS_OA12X4 U908 ( .A(n933), .B(n911), .C(n1036), .Z(
        \mul_b1/result_sat[8] ) );
  HS65_GS_FA1X4 U909 ( .A0(n914), .B0(n913), .CI(n912), .CO(n917), .S0(n915)
         );
  HS65_GS_AO12X4 U910 ( .A(n915), .B(n1036), .C(n933), .Z(
        \mul_b1/result_sat[9] ) );
  HS65_GS_FA1X4 U911 ( .A0(n918), .B0(n917), .CI(n916), .CO(n921), .S0(n919)
         );
  HS65_GS_AO12X4 U912 ( .A(n919), .B(n1036), .C(n933), .Z(
        \mul_b1/result_sat[10] ) );
  HS65_GS_FA1X4 U913 ( .A0(n922), .B0(n921), .CI(n920), .CO(n1032), .S0(n923)
         );
  HS65_GS_OA12X4 U914 ( .A(n933), .B(n923), .C(n1036), .Z(
        \mul_b1/result_sat[11] ) );
  HS65_GSS_XNOR2X3 U915 ( .A(n925), .B(n924), .Z(n927) );
  HS65_GS_OAI21X2 U916 ( .A(n927), .B(n928), .C(n1039), .Z(n926) );
  HS65_GS_CB4I1X4 U917 ( .A(n928), .B(n927), .C(n926), .D(n1036), .Z(
        \mul_b1/result_sat[13] ) );
  HS65_GS_FA1X4 U918 ( .A0(n931), .B0(n930), .CI(n929), .CO(n557), .S0(n932)
         );
  HS65_GS_OA12X4 U919 ( .A(n933), .B(n932), .C(n1036), .Z(
        \mul_b1/result_sat[14] ) );
  HS65_GS_HA1X4 U920 ( .A0(n1020), .B0(n934), .CO(n935), .S0(n963) );
  HS65_GS_PAO2X4 U921 ( .A(\mul_b1/fa1_s1[7] ), .B(n963), .P(x_z2[1]), .Z(
        \mul_b1/fa1_c0[4] ) );
  HS65_GS_HA1X4 U922 ( .A0(n1021), .B0(n935), .CO(n937), .S0(n965) );
  HS65_GS_HA1X4 U923 ( .A0(n1017), .B0(n1016), .CO(n936), .S0(n964) );
  HS65_GS_PAO2X4 U924 ( .A(n965), .B(n964), .P(x_z2[2]), .Z(\mul_b1/fa1_c0[5] ) );
  HS65_GS_HA1X4 U925 ( .A0(n1018), .B0(n936), .CO(n939), .S0(n967) );
  HS65_GS_HA1X4 U926 ( .A0(n1022), .B0(n937), .CO(n938), .S0(n966) );
  HS65_GS_PAO2X4 U927 ( .A(n967), .B(n966), .P(x_z2[3]), .Z(\mul_b1/fa1_c0[6] ) );
  HS65_GS_HA1X4 U928 ( .A0(n1023), .B0(n938), .CO(n940), .S0(n969) );
  HS65_GS_HA1X4 U929 ( .A0(n1019), .B0(n939), .CO(n941), .S0(n968) );
  HS65_GS_PAO2X4 U930 ( .A(n969), .B(n968), .P(x_z2[4]), .Z(\mul_b1/fa1_c0[7] ) );
  HS65_GS_HA1X4 U931 ( .A0(n950), .B0(n940), .CO(n943), .S0(n971) );
  HS65_GS_HA1X4 U932 ( .A0(n1020), .B0(n941), .CO(n942), .S0(n970) );
  HS65_GS_PAO2X4 U933 ( .A(n971), .B(n970), .P(x_z2[5]), .Z(\mul_b1/fa1_c0[8] ) );
  HS65_GS_HA1X4 U934 ( .A0(n1021), .B0(n942), .CO(n944), .S0(n973) );
  HS65_GS_HA1X4 U935 ( .A0(n1024), .B0(n943), .CO(n945), .S0(n972) );
  HS65_GS_PAO2X4 U936 ( .A(n973), .B(n972), .P(x_z2[6]), .Z(\mul_b1/fa1_c0[9] ) );
  HS65_GS_HA1X4 U937 ( .A0(n1022), .B0(n944), .CO(n946), .S0(n975) );
  HS65_GS_HA1X4 U938 ( .A0(n1025), .B0(n945), .CO(n947), .S0(n974) );
  HS65_GS_PAO2X4 U939 ( .A(n975), .B(n974), .P(x_z2[7]), .Z(
        \mul_b1/fa1_c0[10] ) );
  HS65_GS_HA1X4 U940 ( .A0(n1023), .B0(n946), .CO(n949), .S0(n977) );
  HS65_GS_HA1X4 U941 ( .A0(n1026), .B0(n947), .CO(n948), .S0(n976) );
  HS65_GS_PAO2X4 U942 ( .A(n977), .B(n976), .P(x_z2[8]), .Z(
        \mul_b1/fa1_c0[11] ) );
  HS65_GS_HA1X4 U943 ( .A0(n1027), .B0(n948), .CO(n951), .S0(n979) );
  HS65_GS_HA1X4 U944 ( .A0(n950), .B0(n949), .CO(n952), .S0(n978) );
  HS65_GS_PAO2X4 U945 ( .A(n979), .B(n978), .P(x_z2[9]), .Z(
        \mul_b1/fa1_c0[12] ) );
  HS65_GS_HA1X4 U946 ( .A0(n1028), .B0(n951), .CO(n954), .S0(n981) );
  HS65_GS_HA1X4 U947 ( .A0(n1024), .B0(n952), .CO(n953), .S0(n980) );
  HS65_GS_PAO2X4 U948 ( .A(n981), .B(n980), .P(x_z2[10]), .Z(
        \mul_b1/fa1_c0[13] ) );
  HS65_GS_HA1X4 U949 ( .A0(n1025), .B0(n953), .CO(n955), .S0(n983) );
  HS65_GS_HA1X4 U950 ( .A0(n1029), .B0(n954), .CO(n956), .S0(n982) );
  HS65_GS_PAO2X4 U951 ( .A(n983), .B(n982), .P(x_z2[11]), .Z(
        \mul_b1/fa1_c0[14] ) );
  HS65_GS_HA1X4 U952 ( .A0(n1026), .B0(n955), .CO(n958), .S0(n985) );
  HS65_GS_HA1X4 U953 ( .A0(n1030), .B0(n956), .CO(n957), .S0(n984) );
  HS65_GS_PAO2X4 U954 ( .A(n985), .B(n984), .P(x_z2[12]), .Z(
        \mul_b1/fa1_c0[15] ) );
  HS65_GSS_XNOR2X3 U955 ( .A(x_z2[15]), .B(n957), .Z(n987) );
  HS65_GS_HA1X4 U956 ( .A0(n1027), .B0(n958), .CO(n959), .S0(n986) );
  HS65_GS_PAO2X4 U957 ( .A(n987), .B(n986), .P(x_z2[13]), .Z(
        \mul_b1/fa1_c0[16] ) );
  HS65_GS_IVX2 U958 ( .A(n1051), .Z(n962) );
  HS65_GS_HA1X4 U959 ( .A0(n1028), .B0(n959), .CO(n579), .S0(n988) );
  HS65_GS_IVX2 U960 ( .A(n988), .Z(n961) );
  HS65_GS_OAI21X2 U961 ( .A(n1051), .B(n988), .C(x_z2[14]), .Z(n960) );
  HS65_GS_OAI21X2 U962 ( .A(n962), .B(n961), .C(n960), .Z(\mul_b1/fa1_c0[17] )
         );
  HS65_GSS_XOR3X2 U963 ( .A(x_z2[1]), .B(\mul_b1/fa1_s1[7] ), .C(n963), .Z(
        \mul_b1/fa1_s0[4] ) );
  HS65_GSS_XOR3X2 U964 ( .A(x_z2[2]), .B(n965), .C(n964), .Z(
        \mul_b1/fa1_s0[5] ) );
  HS65_GSS_XOR3X2 U965 ( .A(x_z2[3]), .B(n967), .C(n966), .Z(
        \mul_b1/fa1_s0[6] ) );
  HS65_GSS_XOR3X2 U966 ( .A(x_z2[4]), .B(n969), .C(n968), .Z(
        \mul_b1/fa1_s0[7] ) );
  HS65_GSS_XOR3X2 U967 ( .A(x_z2[5]), .B(n971), .C(n970), .Z(
        \mul_b1/fa1_s0[8] ) );
  HS65_GSS_XOR3X2 U968 ( .A(x_z2[6]), .B(n973), .C(n972), .Z(
        \mul_b1/fa1_s0[9] ) );
  HS65_GSS_XOR3X2 U969 ( .A(x_z2[7]), .B(n975), .C(n974), .Z(
        \mul_b1/fa1_s0[10] ) );
  HS65_GSS_XOR3X2 U970 ( .A(x_z2[8]), .B(n977), .C(n976), .Z(
        \mul_b1/fa1_s0[11] ) );
  HS65_GSS_XOR3X2 U971 ( .A(x_z2[9]), .B(n979), .C(n978), .Z(
        \mul_b1/fa1_s0[12] ) );
  HS65_GSS_XOR3X2 U972 ( .A(x_z2[10]), .B(n981), .C(n980), .Z(
        \mul_b1/fa1_s0[13] ) );
  HS65_GSS_XOR3X2 U973 ( .A(x_z2[11]), .B(n983), .C(n982), .Z(
        \mul_b1/fa1_s0[14] ) );
  HS65_GSS_XOR3X2 U974 ( .A(x_z2[12]), .B(n985), .C(n984), .Z(
        \mul_b1/fa1_s0[15] ) );
  HS65_GSS_XOR3X2 U975 ( .A(n987), .B(x_z2[13]), .C(n986), .Z(
        \mul_b1/fa1_s0[16] ) );
  HS65_GSS_XOR3X2 U976 ( .A(n1051), .B(x_z2[14]), .C(n988), .Z(
        \mul_b1/fa1_s0[17] ) );
  HS65_GSS_XNOR2X3 U977 ( .A(n1051), .B(n1030), .Z(n995) );
  HS65_GSS_XNOR2X3 U978 ( .A(n995), .B(n989), .Z(\mul_b1/fa1_s0[18] ) );
  HS65_GSS_XNOR2X3 U979 ( .A(n995), .B(n990), .Z(\mul_b1/fa1_s0[19] ) );
  HS65_GS_HA1X4 U980 ( .A0(n1030), .B0(n991), .CO(n993), .S0(n580) );
  HS65_GSS_XOR2X3 U981 ( .A(x_z2[15]), .B(n993), .Z(n992) );
  HS65_GSS_XNOR2X3 U982 ( .A(n995), .B(n992), .Z(\mul_b1/fa1_s0[20] ) );
  HS65_GS_OR2X4 U983 ( .A(x_z2[15]), .B(n993), .Z(n994) );
  HS65_GSS_XNOR2X3 U984 ( .A(n995), .B(n994), .Z(\mul_b1/fa1_s0[29] ) );
  HS65_GS_MUX21X4 U985 ( .D0(y_z1[5]), .D1(data_out[5]), .S0(valid_in), .Z(
        n3385) );
  HS65_GS_FA1X4 U986 ( .A0(p_a1[4]), .B0(n997), .CI(n996), .CO(n1003), .S0(
        n999) );
  HS65_GS_AOI12X2 U987 ( .A(data_out[4]), .B(n1006), .C(n1005), .Z(n998) );
  HS65_GS_OAI21X2 U988 ( .A(n999), .B(n1008), .C(n998), .Z(n3383) );
  HS65_GS_MUX21X4 U989 ( .D0(y_z1[4]), .D1(data_out[4]), .S0(valid_in), .Z(
        n3382) );
  HS65_GS_MUX21X4 U990 ( .D0(y_z1[3]), .D1(data_out[3]), .S0(valid_in), .Z(
        n3379) );
  HS65_GS_MUX21X4 U991 ( .D0(y_z1[2]), .D1(data_out[2]), .S0(valid_in), .Z(
        n3376) );
  HS65_GS_MUX21X4 U992 ( .D0(y_z1[1]), .D1(data_out[1]), .S0(valid_in), .Z(
        n3373) );
  HS65_GS_CBI4I6X2 U993 ( .A(p_a1[0]), .B(n1001), .C(n1000), .D(n1008), .Z(
        n1002) );
  HS65_GS_AO112X4 U994 ( .A(data_out[0]), .B(n1006), .C(n1002), .D(n1005), .Z(
        n3371) );
  HS65_GS_MUX21X4 U995 ( .D0(\mul_a1/fa1_s2[13] ), .D1(data_out[0]), .S0(
        valid_in), .Z(n3370) );
  HS65_GS_FA1X4 U996 ( .A0(p_a1[5]), .B0(n1004), .CI(n1003), .CO(n785), .S0(
        n1009) );
  HS65_GS_AOI12X2 U997 ( .A(data_out[5]), .B(n1006), .C(n1005), .Z(n1007) );
  HS65_GS_OAI21X2 U998 ( .A(n1009), .B(n1008), .C(n1007), .Z(n3386) );
  HS65_GS_AND2X4 U999 ( .A(\mul_a1/fa1_s2[13] ), .B(n1010), .Z(n1049) );
  HS65_GS_AND2X4 U1000 ( .A(y_z1[1]), .B(n1011), .Z(n1050) );
  HS65_GS_HA1X4 U1001 ( .A0(n1019), .B0(n1012), .CO(n934), .S0(n1013) );
  HS65_GS_AND2X4 U1002 ( .A(\mul_b1/fa1_s1[7] ), .B(n1013), .Z(n1053) );
  HS65_GS_HA1X4 U1003 ( .A0(n1015), .B0(n1014), .CO(n467), .S0(
        \mul_a1/fa1_s1[7] ) );
  HS65_GS_AOI12X2 U1004 ( .A(n1016), .B(n1017), .C(\mul_b1/fa1_c1[8] ), .Z(
        \mul_b1/fa1_s1[8] ) );
  HS65_GS_AOI12X2 U1005 ( .A(n1017), .B(n1018), .C(\mul_b1/fa1_c1[9] ), .Z(
        \mul_b1/fa1_s1[9] ) );
  HS65_GS_AOI12X2 U1006 ( .A(n1018), .B(n1019), .C(\mul_b1/fa1_c1[10] ), .Z(
        \mul_b1/fa1_s1[10] ) );
  HS65_GS_AOI12X2 U1007 ( .A(n1019), .B(n1020), .C(\mul_b1/fa1_c1[11] ), .Z(
        \mul_b1/fa1_s1[11] ) );
  HS65_GS_AOI12X2 U1008 ( .A(n1020), .B(n1021), .C(\mul_b1/fa1_c1[12] ), .Z(
        \mul_b1/fa1_s1[12] ) );
  HS65_GS_AOI12X2 U1009 ( .A(n1021), .B(n1022), .C(\mul_b1/fa1_c1[13] ), .Z(
        \mul_b1/fa1_s1[13] ) );
  HS65_GS_AOI12X2 U1010 ( .A(n1022), .B(n1023), .C(\mul_b1/fa1_c1[14] ), .Z(
        \mul_b1/fa1_s1[14] ) );
  HS65_GS_AOI12X2 U1011 ( .A(n1023), .B(n950), .C(\mul_b1/fa1_c1[15] ), .Z(
        \mul_b1/fa1_s1[15] ) );
  HS65_GS_AOI12X2 U1012 ( .A(n950), .B(n1024), .C(\mul_b1/fa1_c1[16] ), .Z(
        \mul_b1/fa1_s1[16] ) );
  HS65_GS_AOI12X2 U1013 ( .A(n1024), .B(n1025), .C(\mul_b1/fa1_c1[17] ), .Z(
        \mul_b1/fa1_s1[17] ) );
  HS65_GS_AOI12X2 U1014 ( .A(n1025), .B(n1026), .C(\mul_b1/fa1_c1[18] ), .Z(
        \mul_b1/fa1_s1[18] ) );
  HS65_GS_AOI12X2 U1015 ( .A(n1026), .B(n1027), .C(\mul_b1/fa1_c1[19] ), .Z(
        \mul_b1/fa1_s1[19] ) );
  HS65_GS_AOI12X2 U1016 ( .A(n1027), .B(n1028), .C(\mul_b1/fa1_c1[20] ), .Z(
        \mul_b1/fa1_s1[20] ) );
  HS65_GS_AOI12X2 U1017 ( .A(n1028), .B(n1029), .C(\mul_b1/fa1_c1[21] ), .Z(
        \mul_b1/fa1_s1[21] ) );
  HS65_GS_AOI12X2 U1018 ( .A(n1030), .B(n1029), .C(\mul_b1/fa1_c1[22] ), .Z(
        \mul_b1/fa1_s1[22] ) );
  HS65_GS_NOR2X2 U1019 ( .A(n1032), .B(n1033), .Z(n1031) );
  HS65_GS_AOI12X2 U1020 ( .A(n1033), .B(n1032), .C(n1031), .Z(n1034) );
  HS65_GSS_XNOR2X3 U1021 ( .A(n1035), .B(n1034), .Z(n1038) );
  HS65_GS_IVX2 U1022 ( .A(n1036), .Z(n1037) );
  HS65_GS_AOI12X2 U1023 ( .A(n1039), .B(n1038), .C(n1037), .Z(
        \mul_b1/result_sat[12] ) );
  HS65_GS_IVX2 U1024 ( .A(n1040), .Z(n1043) );
  HS65_GS_AOI22X1 U1025 ( .A(n1044), .B(n1043), .C(n1042), .D(n1041), .Z(n1048) );
  HS65_GS_IVX2 U1026 ( .A(n1045), .Z(n1046) );
  HS65_GS_AOI12X2 U1027 ( .A(n1048), .B(n1047), .C(n1046), .Z(
        \mul_b0/result_sat[1] ) );
endmodule

