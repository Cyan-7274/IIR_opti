// 固定系数模块（Q2.14格式、已按matlab排序，最后一节包含总增益）
module opti_coeffs_fixed (
    input  wire [2:0]  stage_index,    // SOS阶段索引(0-5)
    output reg  [15:0] b0,             // 前馈系数b0
    output reg  [15:0] b1,             // 前馈系数b1
    output reg  [15:0] b2,             // 前馈系数b2
    output reg  [15:0] a1,             // 反馈系数a1
    output reg  [15:0] a2              // 反馈系数a2
);
    always @(*) begin
        case (stage_index)
            // 节点1 (原始6)
            3'd0: begin
                b0 = 16'sh4000; // 1.00000000
                b1 = -16'sh2425; // -1.13073730
                b2 = 16'sh4000; // 1.00000000
                a1 = 16'sh4000; // 1.00000000
                a2 = -16'sh3DEF; // -0.96386719
            end
            // 节点2 (原始5)
            3'd1: begin
                b0 = 16'sh4000; // 1.00000000
                b1 = 16'sh2425; // 1.13073730
                b2 = 16'sh4000; // 1.00000000
                a1 = 16'sh4000; // 1.00000000
                a2 = 16'sh3DEF; // 0.96386719
            end
            // 节点3 (原始4)
            3'd2: begin
                b0 = 16'sh4000; // 1.00000000
                b1 = 16'sh294E; // 1.28454590
                b2 = 16'sh4000; // 1.00000000
                a1 = 16'sh4000; // 1.00000000
                a2 = 16'sh332C; // 0.79968262
            end
            // 节点4 (原始3)
            3'd3: begin
                b0 = 16'sh4000; // 1.00000000
                b1 = -16'sh294E; // -1.28454590
                b2 = 16'sh4000; // 1.00000000
                a1 = 16'sh4000; // 1.00000000
                a2 = -16'sh332C; // -0.79968262
            end
            // 节点5 (原始2)
            3'd4: begin
                b0 = 16'sh4000; // 1.00000000
                b1 = -16'sh3950; // -1.79168701
                b2 = 16'sh4000; // 1.00000000
                a1 = 16'sh4000; // 1.00000000
                a2 = -16'sh08E3; // -0.34698486
            end
            // 节点6 (原始1, 含增益)
            3'd5: begin
                b0 = 16'sh01A6; // 0.01544189
                b1 = 16'sh0384; // 0.02770996
                b2 = 16'sh01A6; // 0.01544189
                a1 = 16'sh01A6; // 0.01544189
                a2 = 16'sh0057; // 0.00537109
            end
            default: begin
                b0 = 16'sh4000; b1 = 16'sh0000; b2 = 16'sh0000;
                a1 = 16'sh0000; a2 = 16'sh0000;
            end
        endcase
    end
endmodule